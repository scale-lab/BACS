module buttfly(in_0, in_1, res_0, res_1);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire \add_23/U1.O ;
  wire \add_23/U10.O ;
  wire \add_23/U101.I1 ;
  wire \add_23/U102.I ;
  wire \add_23/U103.I1 ;
  wire \add_23/U104.I ;
  wire \add_23/U105.O ;
  wire \add_23/U112.I1 ;
  wire \add_23/U114.I1 ;
  wire \add_23/U116.I1 ;
  wire \add_23/U117.I ;
  wire \add_23/U118.I1 ;
  wire \add_23/U119.I ;
  wire \add_23/U120.O ;
  wire \add_23/U127.I1 ;
  wire \add_23/U129.I1 ;
  wire \add_23/U131.I1 ;
  wire \add_23/U132.I ;
  wire \add_23/U133.I1 ;
  wire \add_23/U134.I ;
  wire \add_23/U135.O ;
  wire \add_23/U142.I1 ;
  wire \add_23/U144.I1 ;
  wire \add_23/U146.I1 ;
  wire \add_23/U147.I ;
  wire \add_23/U148.I1 ;
  wire \add_23/U149.I ;
  wire \add_23/U150.O ;
  wire \add_23/U157.I1 ;
  wire \add_23/U159.I1 ;
  wire \add_23/U16.I1 ;
  wire \add_23/U161.I1 ;
  wire \add_23/U162.I ;
  wire \add_23/U163.I1 ;
  wire \add_23/U164.I ;
  wire \add_23/U165.O ;
  wire \add_23/U17.I1 ;
  wire \add_23/U172.I1 ;
  wire \add_23/U174.I ;
  wire \add_23/U176.I1 ;
  wire \add_23/U178.I1 ;
  wire \add_23/U18.I ;
  wire \add_23/U180.I ;
  wire \add_23/U182.I1 ;
  wire \add_23/U184.I1 ;
  wire \add_23/U186.I ;
  wire \add_23/U188.I1 ;
  wire \add_23/U19.O ;
  wire \add_23/U190.I1 ;
  wire \add_23/U192.I ;
  wire \add_23/U194.I1 ;
  wire \add_23/U196.I1 ;
  wire \add_23/U198.I ;
  wire \add_23/U200.I1 ;
  wire \add_23/U202.I1 ;
  wire \add_23/U204.I ;
  wire \add_23/U206.I1 ;
  wire \add_23/U208.I1 ;
  wire \add_23/U210.I ;
  wire \add_23/U212.I1 ;
  wire \add_23/U214.I1 ;
  wire \add_23/U216.I ;
  wire \add_23/U218.I1 ;
  wire \add_23/U220.I1 ;
  wire \add_23/U222.I ;
  wire \add_23/U223.I1 ;
  wire \add_23/U225.I1 ;
  wire \add_23/U225.I2 ;
  wire \add_23/U227.I1 ;
  wire \add_23/U228.I ;
  wire \add_23/U229.I1 ;
  wire \add_23/U230.I ;
  wire \add_23/U231.O ;
  wire \add_23/U232.I1 ;
  wire \add_23/U233.I ;
  wire \add_23/U234.I1 ;
  wire \add_23/U235.I ;
  wire \add_23/U25.I1 ;
  wire \add_23/U26.I1 ;
  wire \add_23/U27.I ;
  wire \add_23/U28.O ;
  wire \add_23/U34.I1 ;
  wire \add_23/U35.I1 ;
  wire \add_23/U36.I ;
  wire \add_23/U37.O ;
  wire \add_23/U43.I1 ;
  wire \add_23/U44.I1 ;
  wire \add_23/U45.I ;
  wire \add_23/U46.O ;
  wire \add_23/U52.I1 ;
  wire \add_23/U53.I1 ;
  wire \add_23/U54.I ;
  wire \add_23/U55.O ;
  wire \add_23/U61.I1 ;
  wire \add_23/U62.I1 ;
  wire \add_23/U63.I ;
  wire \add_23/U64.O ;
  wire \add_23/U7.I1 ;
  wire \add_23/U70.I1 ;
  wire \add_23/U71.I1 ;
  wire \add_23/U72.I ;
  wire \add_23/U73.O ;
  wire \add_23/U78.I1 ;
  wire \add_23/U79.I1 ;
  wire \add_23/U8.I1 ;
  wire \add_23/U80.I ;
  wire \add_23/U81.O ;
  wire \add_23/U87.I1 ;
  wire \add_23/U89.I1 ;
  wire \add_23/U9.I ;
  wire \add_23/U90.O ;
  wire \add_23/U97.I1 ;
  wire \add_23/U99.I1 ;
  input [15:0] in_0;
  input [15:0] in_1;
  output [16:0] res_0;
  output [16:0] res_1;
  wire \sub_24/U1.O ;
  wire \sub_24/U100.O ;
  wire \sub_24/U108.I1 ;
  wire \sub_24/U110.I1 ;
  wire \sub_24/U111.I ;
  wire \sub_24/U112.I1 ;
  wire \sub_24/U113.I ;
  wire \sub_24/U114.O ;
  wire \sub_24/U122.I1 ;
  wire \sub_24/U124.I1 ;
  wire \sub_24/U125.I ;
  wire \sub_24/U126.I1 ;
  wire \sub_24/U127.I ;
  wire \sub_24/U128.O ;
  wire \sub_24/U13.I1 ;
  wire \sub_24/U136.I1 ;
  wire \sub_24/U138.I1 ;
  wire \sub_24/U139.I ;
  wire \sub_24/U14.I1 ;
  wire \sub_24/U140.I1 ;
  wire \sub_24/U141.I ;
  wire \sub_24/U142.O ;
  wire \sub_24/U149.I ;
  wire \sub_24/U15.O ;
  wire \sub_24/U151.I ;
  wire \sub_24/U153.I1 ;
  wire \sub_24/U156.I ;
  wire \sub_24/U158.I ;
  wire \sub_24/U160.I1 ;
  wire \sub_24/U163.I ;
  wire \sub_24/U165.I ;
  wire \sub_24/U167.I1 ;
  wire \sub_24/U170.I ;
  wire \sub_24/U172.I ;
  wire \sub_24/U174.I1 ;
  wire \sub_24/U177.I ;
  wire \sub_24/U179.I ;
  wire \sub_24/U181.I1 ;
  wire \sub_24/U184.I ;
  wire \sub_24/U186.I ;
  wire \sub_24/U188.I1 ;
  wire \sub_24/U191.I ;
  wire \sub_24/U193.I ;
  wire \sub_24/U195.I1 ;
  wire \sub_24/U198.I ;
  wire \sub_24/U20.I1 ;
  wire \sub_24/U200.I ;
  wire \sub_24/U202.I1 ;
  wire \sub_24/U205.I ;
  wire \sub_24/U207.I ;
  wire \sub_24/U208.I1 ;
  wire \sub_24/U21.I1 ;
  wire \sub_24/U210.I1 ;
  wire \sub_24/U211.I ;
  wire \sub_24/U212.I1 ;
  wire \sub_24/U213.I ;
  wire \sub_24/U214.O ;
  wire \sub_24/U215.I1 ;
  wire \sub_24/U217.I2 ;
  wire \sub_24/U218.I ;
  wire \sub_24/U22.O ;
  wire \sub_24/U27.I1 ;
  wire \sub_24/U28.I1 ;
  wire \sub_24/U29.O ;
  wire \sub_24/U34.I1 ;
  wire \sub_24/U35.I1 ;
  wire \sub_24/U36.O ;
  wire \sub_24/U41.I1 ;
  wire \sub_24/U42.I1 ;
  wire \sub_24/U43.O ;
  wire \sub_24/U48.I1 ;
  wire \sub_24/U49.I1 ;
  wire \sub_24/U50.O ;
  wire \sub_24/U55.I1 ;
  wire \sub_24/U56.I1 ;
  wire \sub_24/U57.O ;
  wire \sub_24/U6.I1 ;
  wire \sub_24/U62.I1 ;
  wire \sub_24/U63.I1 ;
  wire \sub_24/U64.O ;
  wire \sub_24/U7.I1 ;
  wire \sub_24/U71.I1 ;
  wire \sub_24/U72.O ;
  wire \sub_24/U8.O ;
  wire \sub_24/U80.I1 ;
  wire \sub_24/U82.I1 ;
  wire \sub_24/U83.I ;
  wire \sub_24/U84.I1 ;
  wire \sub_24/U85.I ;
  wire \sub_24/U86.O ;
  wire \sub_24/U94.I1 ;
  wire \sub_24/U96.I1 ;
  wire \sub_24/U97.I ;
  wire \sub_24/U98.I1 ;
  wire \sub_24/U99.I ;
  assign _090_ = ~(in_0[10] ^ in_1[10]);
  assign _091_ = in_1[0] & ~(in_0[0]);
  assign _092_ = in_0[1] & ~(_091_);
  assign _093_ = ~in_0[1];
  assign _094_ = ~((_091_ & _093_) | in_1[1]);
  assign _095_ = ~(_094_ | _092_);
  assign _096_ = in_0[2] & ~(_095_);
  assign _097_ = ~in_0[2];
  assign _098_ = ~((_095_ & _097_) | in_1[2]);
  assign _099_ = ~(_098_ | _096_);
  assign _100_ = in_0[3] & ~(_099_);
  assign _101_ = ~in_0[3];
  assign _102_ = ~((_099_ & _101_) | in_1[3]);
  assign _103_ = ~(_102_ | _100_);
  assign _104_ = in_0[4] & ~(_103_);
  assign _105_ = ~in_0[4];
  assign _106_ = ~((_103_ & _105_) | in_1[4]);
  assign _107_ = ~(_106_ | _104_);
  assign _108_ = in_0[5] & ~(_107_);
  assign _109_ = ~in_0[5];
  assign _110_ = ~((_107_ & _109_) | in_1[5]);
  assign _111_ = ~(_110_ | _108_);
  assign _112_ = in_0[6] & ~(_111_);
  assign _113_ = ~in_0[6];
  assign _114_ = ~((_111_ & _113_) | in_1[6]);
  assign _115_ = ~(_114_ | _112_);
  assign _116_ = in_0[7] & ~(_115_);
  assign _117_ = ~in_0[7];
  assign _118_ = ~((_115_ & _117_) | in_1[7]);
  assign _119_ = ~(_118_ | _116_);
  assign _120_ = in_0[8] & ~(_119_);
  assign _121_ = ~in_0[8];
  assign _122_ = ~((_119_ & _121_) | in_1[8]);
  assign _000_ = ~(_122_ | _120_);
  assign _001_ = in_0[9] & ~(_000_);
  assign _002_ = ~in_0[9];
  assign _003_ = ~((_000_ & _002_) | in_1[9]);
  assign _004_ = ~(_003_ | _001_);
  assign \sub_24/U142.O  = ~(_004_ ^ _090_);
  assign _005_ = ~(in_0[11] ^ in_1[11]);
  assign _006_ = in_0[10] & ~(_004_);
  assign _007_ = ~in_0[10];
  assign _008_ = ~((_004_ & _007_) | in_1[10]);
  assign _009_ = ~(_008_ | _006_);
  assign \sub_24/U128.O  = ~(_009_ ^ _005_);
  assign _010_ = ~(in_0[12] ^ in_1[12]);
  assign _011_ = in_0[11] & ~(_009_);
  assign _012_ = ~in_0[11];
  assign _013_ = ~((_009_ & _012_) | in_1[11]);
  assign _014_ = ~(_013_ | _011_);
  assign \sub_24/U114.O  = ~(_014_ ^ _010_);
  assign _015_ = ~(in_0[13] ^ in_1[13]);
  assign _016_ = in_0[12] & ~(_014_);
  assign _017_ = ~in_0[12];
  assign _018_ = ~((_014_ & _017_) | in_1[12]);
  assign _019_ = ~(_018_ | _016_);
  assign \sub_24/U100.O  = ~(_019_ ^ _015_);
  assign _020_ = ~(in_0[14] ^ in_1[14]);
  assign _021_ = in_0[13] & ~(_019_);
  assign _022_ = ~in_0[13];
  assign _023_ = ~((_019_ & _022_) | in_1[13]);
  assign _024_ = ~(_023_ | _021_);
  assign \sub_24/U86.O  = ~(_024_ ^ _020_);
  assign _025_ = ~(in_0[15] ^ in_1[15]);
  assign _026_ = ~_025_;
  assign _027_ = in_0[14] & ~(_024_);
  assign _028_ = ~in_0[14];
  assign _029_ = ~((_024_ & _028_) | in_1[14]);
  assign _030_ = ~(_029_ | _027_);
  assign \sub_24/U72.O  = _030_ ^ _026_;
  assign _031_ = ~in_0[15];
  assign _032_ = _030_ | _031_;
  assign _033_ = ~((_030_ & _031_) | in_1[15]);
  assign _034_ = _032_ & ~(_033_);
  assign \sub_24/U64.O  = _034_ ^ _026_;
  assign _035_ = ~(in_1[1] ^ in_0[1]);
  assign \sub_24/U57.O  = ~(_035_ ^ _091_);
  assign _036_ = ~(in_1[2] ^ in_0[2]);
  assign \sub_24/U50.O  = ~(_036_ ^ _095_);
  assign _037_ = ~(in_1[3] ^ in_0[3]);
  assign \sub_24/U43.O  = ~(_037_ ^ _099_);
  assign _038_ = ~(in_1[4] ^ in_0[4]);
  assign \sub_24/U36.O  = ~(_038_ ^ _103_);
  assign _039_ = ~(in_1[5] ^ in_0[5]);
  assign \sub_24/U29.O  = ~(_039_ ^ _107_);
  assign _040_ = ~(in_1[6] ^ in_0[6]);
  assign \sub_24/U22.O  = ~(_040_ ^ _111_);
  assign _041_ = ~(in_1[7] ^ in_0[7]);
  assign \sub_24/U15.O  = ~(_041_ ^ _115_);
  assign _042_ = ~(in_1[8] ^ in_0[8]);
  assign \sub_24/U8.O  = ~(_042_ ^ _119_);
  assign _043_ = ~(in_1[9] ^ in_0[9]);
  assign \sub_24/U1.O  = ~(_043_ ^ _000_);
  assign \add_23/U231.O  = in_0[0] ^ in_1[0];
  assign _044_ = ~(in_0[0] & in_1[0]);
  assign \add_23/U73.O  = _044_ ^ _035_;
  assign _045_ = in_0[1] & ~(_044_);
  assign _046_ = ~(_044_ & _093_);
  assign _047_ = ~((_046_ & in_1[1]) | _045_);
  assign _048_ = in_0[2] & ~(_047_);
  assign _049_ = ~(_047_ & _097_);
  assign _050_ = ~((_049_ & in_1[2]) | _048_);
  assign _051_ = in_0[3] & ~(_050_);
  assign _052_ = ~(_050_ & _101_);
  assign _053_ = ~((_052_ & in_1[3]) | _051_);
  assign _054_ = in_0[4] & ~(_053_);
  assign _055_ = ~(_053_ & _105_);
  assign _056_ = ~((_055_ & in_1[4]) | _054_);
  assign _057_ = in_0[5] & ~(_056_);
  assign _058_ = ~(_056_ & _109_);
  assign _059_ = ~((_058_ & in_1[5]) | _057_);
  assign _060_ = in_0[6] & ~(_059_);
  assign _061_ = ~(_059_ & _113_);
  assign _062_ = ~((_061_ & in_1[6]) | _060_);
  assign _063_ = in_0[7] & ~(_062_);
  assign _064_ = ~(_062_ & _117_);
  assign _065_ = ~((_064_ & in_1[7]) | _063_);
  assign _066_ = in_0[8] & ~(_065_);
  assign _067_ = ~(_065_ & _121_);
  assign _068_ = ~((_067_ & in_1[8]) | _066_);
  assign _069_ = in_0[9] & ~(_068_);
  assign _070_ = ~(_068_ & _002_);
  assign _071_ = ~((_070_ & in_1[9]) | _069_);
  assign \add_23/U165.O  = _071_ ^ _090_;
  assign _072_ = in_0[10] & ~(_071_);
  assign _073_ = ~(_071_ & _007_);
  assign _074_ = ~((_073_ & in_1[10]) | _072_);
  assign \add_23/U150.O  = _074_ ^ _005_;
  assign _075_ = in_0[11] & ~(_074_);
  assign _076_ = ~(_074_ & _012_);
  assign _077_ = ~((_076_ & in_1[11]) | _075_);
  assign \add_23/U135.O  = _077_ ^ _010_;
  assign _078_ = in_0[12] & ~(_077_);
  assign _079_ = ~(_077_ & _017_);
  assign _080_ = ~((_079_ & in_1[12]) | _078_);
  assign \add_23/U120.O  = _080_ ^ _015_;
  assign _081_ = in_0[13] & ~(_080_);
  assign _082_ = ~(_080_ & _022_);
  assign _083_ = ~((_082_ & in_1[13]) | _081_);
  assign \add_23/U105.O  = _083_ ^ _020_;
  assign _084_ = in_0[14] & ~(_083_);
  assign _085_ = ~(_083_ & _028_);
  assign _086_ = ~((_085_ & in_1[14]) | _084_);
  assign \add_23/U90.O  = _086_ ^ _025_;
  assign _087_ = in_0[15] & ~(_086_);
  assign _088_ = ~(_086_ & _031_);
  assign _089_ = ~((_088_ & in_1[15]) | _087_);
  assign \add_23/U81.O  = _089_ ^ _025_;
  assign \add_23/U64.O  = _047_ ^ _036_;
  assign \add_23/U55.O  = _050_ ^ _037_;
  assign \add_23/U46.O  = _053_ ^ _038_;
  assign \add_23/U37.O  = _056_ ^ _039_;
  assign \add_23/U28.O  = _059_ ^ _040_;
  assign \add_23/U19.O  = _062_ ^ _041_;
  assign \add_23/U10.O  = _065_ ^ _042_;
  assign \add_23/U1.O  = _068_ ^ _043_;
  assign \sub_24/U56.I1  = in_0[2];
  assign \sub_24/U193.I  = in_0[3];
  assign \add_23/U63.I  = in_1[3];
  assign \add_23/U62.I1  = in_0[3];
  assign \add_23/U61.I1  = in_1[3];
  assign \sub_24/U195.I1  = in_0[3];
  assign \sub_24/U6.I1  = in_1[9];
  assign \sub_24/U160.I1  = in_0[8];
  assign \sub_24/U110.I1  = in_1[13];
  assign \sub_24/U62.I1  = in_1[1];
  assign \sub_24/U63.I1  = in_0[1];
  assign \sub_24/U136.I1  = in_0[10];
  assign \add_23/U16.I1  = in_1[8];
  assign \add_23/U144.I1  = in_0[11];
  assign \add_23/U54.I  = in_1[4];
  assign \sub_24/U198.I  = in_1[2];
  assign \add_23/U53.I1  = in_0[4];
  assign \add_23/U52.I1  = in_1[4];
  assign \add_23/U161.I1  = in_1[11];
  assign \sub_24/U163.I  = in_1[7];
  assign \sub_24/U7.I1  = in_0[9];
  assign res_1 = { \sub_24/U64.O , \sub_24/U72.O , \sub_24/U86.O , \sub_24/U100.O , \sub_24/U114.O , \sub_24/U128.O , \sub_24/U142.O , \sub_24/U1.O , \sub_24/U8.O , \sub_24/U15.O , \sub_24/U22.O , \sub_24/U29.O , \sub_24/U36.O , \sub_24/U43.O , \sub_24/U50.O , \sub_24/U57.O , \add_23/U231.O  };
  assign \sub_24/U111.I  = in_0[13];
  assign \sub_24/U138.I1  = in_1[11];
  assign \sub_24/U71.I1  = in_0[15];
  assign \sub_24/U20.I1  = in_1[7];
  assign \sub_24/U165.I  = in_0[7];
  assign \add_23/U162.I  = in_0[11];
  assign \sub_24/U122.I1  = in_0[11];
  assign \sub_24/U200.I  = in_0[2];
  assign \sub_24/U139.I  = in_0[11];
  assign \add_23/U45.I  = in_1[5];
  assign \sub_24/U167.I1  = in_0[7];
  assign \add_23/U163.I1  = in_0[11];
  assign \add_23/U44.I1  = in_0[5];
  assign \sub_24/U202.I1  = in_0[2];
  assign res_0 = { \add_23/U81.O , \add_23/U90.O , \add_23/U105.O , \add_23/U120.O , \add_23/U135.O , \add_23/U150.O , \add_23/U165.O , \add_23/U1.O , \add_23/U10.O , \add_23/U19.O , \add_23/U28.O , \add_23/U37.O , \add_23/U46.O , \add_23/U55.O , \add_23/U64.O , \add_23/U73.O , \add_23/U231.O  };
  assign \add_23/U43.I1  = in_1[5];
  assign \add_23/U164.I  = in_1[11];
  assign \sub_24/U14.I1  = in_0[8];
  assign \sub_24/U80.I1  = in_0[14];
  assign \sub_24/U112.I1  = in_0[13];
  assign \add_23/U118.I1  = in_0[14];
  assign \sub_24/U82.I1  = in_1[15];
  assign \sub_24/U140.I1  = in_0[11];
  assign \sub_24/U83.I  = in_0[15];
  assign \sub_24/U84.I1  = in_0[15];
  assign \sub_24/U205.I  = in_1[1];
  assign \sub_24/U85.I  = in_1[15];
  assign \sub_24/U124.I1  = in_1[12];
  assign \add_23/U36.I  = in_1[6];
  assign \sub_24/U141.I  = in_1[11];
  assign \add_23/U35.I1  = in_0[6];
  assign \sub_24/U113.I  = in_1[13];
  assign \sub_24/U170.I  = in_1[6];
  assign \add_23/U34.I1  = in_1[6];
  assign \sub_24/U207.I  = in_0[1];
  assign \sub_24/U208.I1  = in_0[1];
  assign \sub_24/U172.I  = in_0[6];
  assign \sub_24/U125.I  = in_0[12];
  assign \sub_24/U21.I1  = in_0[7];
  assign \sub_24/U94.I1  = in_0[13];
  assign \add_23/U146.I1  = in_1[12];
  assign \add_23/U27.I  = in_1[7];
  assign \sub_24/U96.I1  = in_1[14];
  assign \sub_24/U97.I  = in_0[14];
  assign \add_23/U26.I1  = in_0[7];
  assign \sub_24/U98.I1  = in_0[14];
  assign \sub_24/U210.I1  = in_1[10];
  assign \sub_24/U174.I1  = in_0[6];
  assign \sub_24/U99.I  = in_1[14];
  assign \add_23/U25.I1  = in_1[7];
  assign \sub_24/U126.I1  = in_0[12];
  assign \sub_24/U211.I  = in_0[10];
  assign \add_23/U235.I  = in_1[0];
  assign \add_23/U234.I1  = in_0[0];
  assign \sub_24/U212.I1  = in_0[10];
  assign \add_23/U233.I  = in_0[0];
  assign \add_23/U232.I1  = in_1[0];
  assign \sub_24/U127.I  = in_1[12];
  assign \add_23/U230.I  = in_1[10];
  assign \sub_24/U213.I  = in_1[10];
  assign \add_23/U99.I1  = in_0[14];
  assign \add_23/U147.I  = in_0[12];
  assign \add_23/U229.I1  = in_0[10];
  assign \sub_24/U214.O  = \add_23/U231.O ;
  assign \add_23/U228.I  = in_0[10];
  assign \sub_24/U215.I1  = in_0[0];
  assign \add_23/U227.I1  = in_1[10];
  assign \add_23/U225.I2  = in_0[0];
  assign \add_23/U225.I1  = in_1[0];
  assign \add_23/U97.I1  = in_1[14];
  assign \sub_24/U177.I  = in_1[5];
  assign \sub_24/U217.I2  = in_0[0];
  assign \add_23/U223.I1  = in_0[1];
  assign \add_23/U222.I  = in_0[1];
  assign \sub_24/U218.I  = in_1[0];
  assign \add_23/U220.I1  = in_1[1];
  assign \add_23/U218.I1  = in_0[2];
  assign \add_23/U216.I  = in_0[2];
  assign \sub_24/U179.I  = in_0[5];
  assign \add_23/U117.I  = in_0[14];
  assign \sub_24/U149.I  = in_1[9];
  assign \add_23/U214.I1  = in_1[2];
  assign \add_23/U148.I1  = in_0[12];
  assign \sub_24/U27.I1  = in_1[6];
  assign \add_23/U212.I1  = in_0[3];
  assign \add_23/U142.I1  = in_1[11];
  assign \add_23/U210.I  = in_0[3];
  assign \sub_24/U28.I1  = in_0[6];
  assign \add_23/U9.I  = in_1[9];
  assign \sub_24/U181.I1  = in_0[5];
  assign \add_23/U116.I1  = in_1[14];
  assign \add_23/U157.I1  = in_1[10];
  assign \add_23/U89.I1  = in_0[15];
  assign \add_23/U208.I1  = in_1[3];
  assign \add_23/U206.I1  = in_0[4];
  assign \add_23/U87.I1  = in_1[15];
  assign \sub_24/U13.I1  = in_1[8];
  assign \add_23/U204.I  = in_0[4];
  assign \add_23/U149.I  = in_1[12];
  assign \sub_24/U151.I  = in_0[9];
  assign \sub_24/U34.I1  = in_1[5];
  assign \add_23/U202.I1  = in_1[4];
  assign \sub_24/U108.I1  = in_0[12];
  assign \add_23/U102.I  = in_0[15];
  assign \sub_24/U35.I1  = in_0[5];
  assign \sub_24/U184.I  = in_1[4];
  assign \add_23/U200.I1  = in_0[5];
  assign \add_23/U198.I  = in_0[5];
  assign \add_23/U80.I  = in_1[1];
  assign \add_23/U114.I1  = in_0[13];
  assign \add_23/U196.I1  = in_1[5];
  assign \add_23/U8.I1  = in_0[9];
  assign \add_23/U134.I  = in_1[13];
  assign \sub_24/U153.I1  = in_0[9];
  assign \add_23/U79.I1  = in_0[1];
  assign \add_23/U194.I1  = in_0[6];
  assign \sub_24/U186.I  = in_0[4];
  assign \add_23/U78.I1  = in_1[1];
  assign \add_23/U192.I  = in_0[6];
  assign \add_23/U133.I1  = in_0[13];
  assign \sub_24/U41.I1  = in_1[4];
  assign \add_23/U132.I  = in_0[13];
  assign \add_23/U190.I1  = in_1[6];
  assign \sub_24/U42.I1  = in_0[4];
  assign \add_23/U119.I  = in_1[14];
  assign \sub_24/U188.I1  = in_0[4];
  assign \add_23/U188.I1  = in_0[7];
  assign \add_23/U131.I1  = in_1[13];
  assign \add_23/U186.I  = in_0[7];
  assign \add_23/U101.I1  = in_1[15];
  assign \add_23/U184.I1  = in_1[7];
  assign \add_23/U182.I1  = in_0[8];
  assign \add_23/U72.I  = in_1[2];
  assign \add_23/U180.I  = in_0[8];
  assign \sub_24/U48.I1  = in_1[3];
  assign \add_23/U18.I  = in_1[8];
  assign \add_23/U71.I1  = in_0[2];
  assign \sub_24/U156.I  = in_1[8];
  assign \sub_24/U49.I1  = in_0[3];
  assign \add_23/U70.I1  = in_1[2];
  assign \add_23/U178.I1  = in_1[8];
  assign \add_23/U129.I1  = in_0[12];
  assign \add_23/U7.I1  = in_1[9];
  assign \add_23/U176.I1  = in_0[9];
  assign \add_23/U159.I1  = in_0[10];
  assign \add_23/U174.I  = in_0[9];
  assign \add_23/U112.I1  = in_1[13];
  assign \sub_24/U191.I  = in_1[3];
  assign \add_23/U172.I1  = in_1[9];
  assign \sub_24/U158.I  = in_0[8];
  assign \add_23/U103.I1  = in_0[15];
  assign \add_23/U127.I1  = in_1[12];
  assign \add_23/U17.I1  = in_0[8];
  assign \sub_24/U55.I1  = in_1[2];
  assign \add_23/U104.I  = in_1[15];
endmodule
