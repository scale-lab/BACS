module sad (a,b,c,d,e,f,out,clk,rst);

input clk, rst;
input [7:0] a,b,c,d,e,f;
output [32:0] out;

wire [7:0] sa,sb,sc,sd,se,sf;
wire [8:0] da,db,dc;
wire [8:0] dadb,dadbdc;
wire [2:0] carry;

wire b0,b1,b2,c0,c1;
wire s0,s1,s2,s3,s4,s5,s6;

reg [31:0] accum;

assign sa=(a>=b)?a:b;
assign sb=(a>=b)?b:a;
assign sc=(c>=d)?c:d;
assign sd=(c>=d)?d:c;
assign se=(e>=f)?e:f;
assign sf=(e>=f)?f:e;

//sub8 U1 (.a(sa),.b(sb),.r(da));
sub4_bin U00 (.in({sb[3:0],sa[3:0],1'b0}),.out({b0,da[3:0]}));
sub4_bin U01 (.in({sb[7:4],sa[7:4],b0}),.out(da[8:4]));
//sub8 U2 (.a(sc),.b(sd),.r(db));
sub4_bin U02 (.in({sd[3:0],sc[3:0],1'b0}),.out({b1,db[3:0]}));
sub4_bin U03 (.in({sd[7:4],sc[7:4],b1}),.out(db[8:4]));
//sub8 U3 (.a(se),.b(sf),.r(dc));
sub4_bin U04 (.in({sf[3:0],se[3:0],1'b0}),.out({b2,dc[3:0]}));
sub4_bin U05 (.in({sf[7:4],se[7:4],b2}),.out(dc[8:4]));

//adder8 U4 (.a(da[7:0]),.b(db[7:0]),.r(dadb));
add4_cin U06 (.in({db[3:0],da[3:0],1'b0}),.out({c0,dadb[3:0]}));
add4_cin U07 (.in({db[7:4],da[7:4],c0}),.out(dadb[8:4]));
//adder8 U5 (.a(dadb[7:0]),.b(dc[7:0]),.r(dadbdc));
add4_cin U08 (.in({b[3:0],a[3:0],1'b0}),.out({c1,dadbdc[3:0]}));
add4_cin U09 (.in({b[7:4],a[7:4],c1}),.out(dadbdc[8:4]));

assign carry=dadb[8]+dadbdc[8]+da[8]+db[8]+dc[8];

//adder32 U6 (.a({21'b0,carry,dadbdc[7:0]}),.b(accum),.r(out));
add4_cin U10 (.in({accum[3:0],dadbdc[3:0],1'b0}),.out({s0,out[3:0]}));
add4_cin U11 (.in({accum[7:4],dadbdc[7:4],s0}),.out({s1,out[7:4]}));
add4_cin U12 (.in({accum[11:8],4'b0000,s1}),.out({s2,out[11:8]}));
add4_cin U13 (.in({accum[15:12],4'b0000,s2}),.out({s3,out[15:12]}));
add4_cin U14 (.in({accum[19:16],4'b0000,s3}),.out({s4,out[19:16]}));
add4_cin U15 (.in({accum[23:20],4'b0000,s4}),.out({s5,out[23:20]}));
add4_cin U16 (.in({accum[27:24],4'b0000,s5}),.out({s6,out[27:24]}));
add4_cin U17 (.in({accum[31:28],4'b0000,s6}),.out(out[32:28]));


always@(posedge clk or negedge rst)
begin
    if(!rst)
        accum<=32'b0;
    else
        accum<=out[31:0];
end

endmodule

module sub4_bin (
input [8:0] in,
output [4:0] out);

assign out[4] = (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]);
assign out[3] = (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]);
assign out[2] = (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]);
assign out[1] = (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]);
assign out[0] = (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]);

endmodule

module add4_cin (
input [8:0] in,
output [4:0] out);

assign out[4] = (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]);
assign out[3] = (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]);
assign out[2] = (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]);
assign out[1] = (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]);
assign out[0] = (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]);

endmodule
