
module add4_cin(
input [8:0] in,
output [4:0] out);

assign out[4] = (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]);
assign out[3] = (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]);
assign out[2] = (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]);
assign out[1] = (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]);
assign out[0] = (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]);

endmodule

