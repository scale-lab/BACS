module sad (a,b,c,d,e,f,out,clk,rst);

input clk, rst;
input [7:0] a,b,c,d,e,f;
output [32:0] out;

wire [7:0] sa,sb,sc,sd,se,sf;
wire [8:0] da,db,dc;
wire [8:0] dadb,dadbdc;
wire [2:0] carry;

reg [31:0] accum;

assign sa=(a>=b)?a:b;
assign sb=(a>=b)?b:a;
assign sc=(c>=d)?c:d;
assign sd=(c>=d)?d:c;
assign se=(e>=f)?e:f;
assign sf=(e>=f)?f:e;

sub8 U1 (.a(sa),.b(sb),.r(da));
sub8 U2 (.a(sc),.b(sd),.r(db));
sub8 U3 (.a(se),.b(sf),.r(dc));

adder8 U4 (.a(da[7:0]),.b(db[7:0]),.r(dadb));
adder8 U5 (.a(dadb[7:0]),.b(dc[7:0]),.r(dadbdc));

assign carry=dadb[8]+dadbdc[8]+da[8]+db[8]+dc[8];

adder32 U6 (.a({21'b0,carry,dadbdc[7:0]}),.b(accum),.r(out));

always@(posedge clk or negedge rst)
begin
    if(!rst)
        accum<=32'b0;
    else
        accum<=out[31:0];
end

endmodule

module sub8 (a,b,r);

input [7:0] a,b;
output [8:0] r;

wire [4:0] s0,s1;

sub4_bin U1 (.in({b[3:0],a[3:0],1'b0}),.out(s0));
sub4_bin U2 (.in({b[7:4],a[7:4],s0[4]}),.out(s1));

assign r={s1,s0[3:0]};

endmodule
module adder8 (a,b,r);

input [7:0] a,b;
output [8:0] r;

wire [4:0] s0,s1;

add4_cin U1 (.in({b[3:0],a[3:0],1'b0}),.out(s0));
add4_cin U2 (.in({b[7:4],a[7:4],s0[4]}),.out(s1));

assign r={s1,s0[3:0]};

endmodule
module adder32 (a,b,r);

input [31:0] a,b;
output [32:0] r;

wire [4:0] s0,s1,s2,s3,s4,s5,s6,s7;

add4_cin U1 (.in({b[3:0],a[3:0],1'b0}),.out(s0));
add4_cin U2 (.in({b[7:4],a[7:4],s0[4]}),.out(s1));
add4_cin U3 (.in({b[11:8],a[11:8],s1[4]}),.out(s2));
add4_cin U4 (.in({b[15:12],a[15:12],s2[4]}),.out(s3));
add4_cin U5 (.in({b[19:16],a[19:16],s3[4]}),.out(s4));
add4_cin U6 (.in({b[23:20],a[23:20],s4[4]}),.out(s5));
add4_cin U7 (.in({b[27:24],a[27:24],s5[4]}),.out(s6));
add4_cin U8 (.in({b[31:28],a[31:28],s6[4]}),.out(s7));

assign r={s7,s6[3:0],s5[3:0],s4[3:0],s3[3:0],s2[3:0],s1[3:0],s0[3:0]};

endmodule
module add4(
input [7:0] in,
output [4:0] out);

assign out[4] = (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7]);
assign out[3] = (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7]);
assign out[2] = (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7]);
assign out[1] = (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7]);
assign out[0] = (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7]);

endmodule
module sub4_bin(
input [8:0] in,
output [4:0] out);

assign out[4] = (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]);
assign out[3] = (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]);
assign out[2] = (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]);
assign out[1] = (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]);
assign out[0] = (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]);

endmodule
