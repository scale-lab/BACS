module but (a,b,sum,diff);

input [7:0] a,b;
output [8:0] sum, diff;

wire c0,b0;
wire [7:0] sa,sb;

assign sa=(a>=b)?a:b;
assign sb=(a>=b)?b:a;

//adder8 U0 (.a(sa),.b(sb),.r(sum));
add4_cin U0 (.in({sa[3:0],sb[3:0],1'b0}),.out({c0,sum[3:0]}));
add4_cin U1 (.in({sa[7:4],sb[7:4],c0}),.out(sum[8:4]));

//sub8 U1 (.a(sa),.b(sb),.r(diff));
sub4_bin U2 (.in({sb[3:0],sa[3:0],1'b0}),.out({b0,diff[3:0]}));
sub4_bin U3 (.in({sb[7:4],sa[7:4],b0}),.out(diff[8:4]));


endmodule

module add4_cin(
input [8:0] in,
output [4:0] out);

assign out[4] = (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]);
assign out[3] = (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]);
assign out[2] = (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]);
assign out[1] = (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]);
assign out[0] = (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]);

endmodule
module sub4_bin(
input [8:0] in,
output [4:0] out);

assign out[4] = (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]);
assign out[3] = (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]);
assign out[2] = (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]);
assign out[1] = (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]);
assign out[0] = (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(~in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(~in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(~in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(~in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(~in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(~in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(~in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (~in[0])&(~in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]) | (in[0])&(in[1])&(in[2])&(in[3])&(in[4])&(in[5])&(in[6])&(in[7])&(in[8]);

endmodule
