module sin_tb;
reg [23:0] pi;
wire [24:0] po;
sin dut( pi[0] , pi[1] , pi[2] , pi[3] , pi[4] , pi[5] , pi[6] , pi[7] , pi[8] , pi[9] , pi[10] , pi[11] , pi[12] , pi[13] , pi[14] , pi[15] , pi[16] , pi[17] , pi[18] , pi[19] , pi[20] , pi[21] , pi[22] , pi[23] , po[0] , po[1] , po[2] , po[3] , po[4] , po[5] , po[6] , po[7] , po[8] , po[9] , po[10] , po[11] , po[12] , po[13] , po[14] , po[15] , po[16] , po[17] , po[18] , po[19] , po[20] , po[21] , po[22] , po[23] , po[24] );
initial
begin
# 1  pi=24'b011101010000010011000010;
#1 $display("%b", po);
# 1  pi=24'b100011011000101010100001;
#1 $display("%b", po);
# 1  pi=24'b100000100111000111101000;
#1 $display("%b", po);
# 1  pi=24'b101110010011011100101010;
#1 $display("%b", po);
# 1  pi=24'b000011000011011000001000;
#1 $display("%b", po);
# 1  pi=24'b100100011011100010011101;
#1 $display("%b", po);
# 1  pi=24'b100010100100101100111110;
#1 $display("%b", po);
# 1  pi=24'b110110001100111100100011;
#1 $display("%b", po);
# 1  pi=24'b001101100011010110011011;
#1 $display("%b", po);
# 1  pi=24'b000001011001001001100110;
#1 $display("%b", po);
# 1  pi=24'b011111001101110000101100;
#1 $display("%b", po);
# 1  pi=24'b110010011101101100000110;
#1 $display("%b", po);
# 1  pi=24'b000100110100011001010010;
#1 $display("%b", po);
# 1  pi=24'b110110101010110111101011;
#1 $display("%b", po);
# 1  pi=24'b001110100101110000100011;
#1 $display("%b", po);
# 1  pi=24'b111000011001011011001111;
#1 $display("%b", po);
# 1  pi=24'b100011110011101000111001;
#1 $display("%b", po);
# 1  pi=24'b111100010010000011110111;
#1 $display("%b", po);
# 1  pi=24'b000001101011011101111100;
#1 $display("%b", po);
# 1  pi=24'b110000000001111001010100;
#1 $display("%b", po);
# 1  pi=24'b110000011100110011110011;
#1 $display("%b", po);
# 1  pi=24'b000010100110001110001001;
#1 $display("%b", po);
# 1  pi=24'b000101001111010011000011;
#1 $display("%b", po);
# 1  pi=24'b100000101110010100110101;
#1 $display("%b", po);
# 1  pi=24'b001011101110001101000010;
#1 $display("%b", po);
# 1  pi=24'b101101000011011010110011;
#1 $display("%b", po);
# 1  pi=24'b111111001011111001010010;
#1 $display("%b", po);
# 1  pi=24'b000110101011100001001111;
#1 $display("%b", po);
# 1  pi=24'b101100101011011100000011;
#1 $display("%b", po);
# 1  pi=24'b111101000000001000111110;
#1 $display("%b", po);
# 1  pi=24'b011100010101110010000010;
#1 $display("%b", po);
# 1  pi=24'b010011001101111011011101;
#1 $display("%b", po);
# 1  pi=24'b010011001101100000111011;
#1 $display("%b", po);
# 1  pi=24'b110010110001011100010001;
#1 $display("%b", po);
# 1  pi=24'b100101001111010101110111;
#1 $display("%b", po);
# 1  pi=24'b110011100010001000111100;
#1 $display("%b", po);
# 1  pi=24'b100111001100010010011101;
#1 $display("%b", po);
# 1  pi=24'b001111011110011000111011;
#1 $display("%b", po);
# 1  pi=24'b011111111001011000110000;
#1 $display("%b", po);
# 1  pi=24'b011101000111010001101010;
#1 $display("%b", po);
# 1  pi=24'b001000000110001001101100;
#1 $display("%b", po);
# 1  pi=24'b000111011000110001111010;
#1 $display("%b", po);
# 1  pi=24'b101001101100000101101100;
#1 $display("%b", po);
# 1  pi=24'b000011101000100111001100;
#1 $display("%b", po);
# 1  pi=24'b000111000010000101101011;
#1 $display("%b", po);
# 1  pi=24'b101101101100010111110111;
#1 $display("%b", po);
# 1  pi=24'b010001110000000000011100;
#1 $display("%b", po);
# 1  pi=24'b001010110101110100000100;
#1 $display("%b", po);
# 1  pi=24'b101011100001001000100000;
#1 $display("%b", po);
# 1  pi=24'b110111110101001011001000;
#1 $display("%b", po);
# 1  pi=24'b110000000110101101101101;
#1 $display("%b", po);
# 1  pi=24'b000101110100011100011110;
#1 $display("%b", po);
# 1  pi=24'b001100110011110110010000;
#1 $display("%b", po);
# 1  pi=24'b101010111100000000100000;
#1 $display("%b", po);
# 1  pi=24'b100010100011110110010000;
#1 $display("%b", po);
# 1  pi=24'b101010110110110101010001;
#1 $display("%b", po);
# 1  pi=24'b111110110100001101100011;
#1 $display("%b", po);
# 1  pi=24'b100100110000100101000111;
#1 $display("%b", po);
# 1  pi=24'b010111010011100010111110;
#1 $display("%b", po);
# 1  pi=24'b110111010101010000101111;
#1 $display("%b", po);
# 1  pi=24'b110101001010010000001100;
#1 $display("%b", po);
# 1  pi=24'b010110010101100110011101;
#1 $display("%b", po);
# 1  pi=24'b011010001010110101011010;
#1 $display("%b", po);
# 1  pi=24'b111111011010110101000000;
#1 $display("%b", po);
# 1  pi=24'b010100000101011000011101;
#1 $display("%b", po);
# 1  pi=24'b000000010101100001001100;
#1 $display("%b", po);
# 1  pi=24'b111011100110010110011011;
#1 $display("%b", po);
# 1  pi=24'b011000010010101000100111;
#1 $display("%b", po);
# 1  pi=24'b101101011101000110001101;
#1 $display("%b", po);
# 1  pi=24'b000011000111001001100111;
#1 $display("%b", po);
# 1  pi=24'b100000111011000110101001;
#1 $display("%b", po);
# 1  pi=24'b000001000111101110100011;
#1 $display("%b", po);
# 1  pi=24'b010010001110111011010101;
#1 $display("%b", po);
# 1  pi=24'b000000001010100111110001;
#1 $display("%b", po);
# 1  pi=24'b111010011111000010000011;
#1 $display("%b", po);
# 1  pi=24'b111111100011101101000011;
#1 $display("%b", po);
# 1  pi=24'b000111100010000101011101;
#1 $display("%b", po);
# 1  pi=24'b100101111001111110100000;
#1 $display("%b", po);
# 1  pi=24'b101001110011010100011011;
#1 $display("%b", po);
# 1  pi=24'b111111100110011011110100;
#1 $display("%b", po);
# 1  pi=24'b000111110101110111110000;
#1 $display("%b", po);
# 1  pi=24'b110101111000011101000000;
#1 $display("%b", po);
# 1  pi=24'b011111110010010000001011;
#1 $display("%b", po);
# 1  pi=24'b101010111011001001011000;
#1 $display("%b", po);
# 1  pi=24'b110100101011110110101010;
#1 $display("%b", po);
# 1  pi=24'b000110101101000001111000;
#1 $display("%b", po);
# 1  pi=24'b100111011011001011100010;
#1 $display("%b", po);
# 1  pi=24'b000000001111110101101111;
#1 $display("%b", po);
# 1  pi=24'b011110101000000010001101;
#1 $display("%b", po);
# 1  pi=24'b110010101100110100000011;
#1 $display("%b", po);
# 1  pi=24'b110101000011011000001101;
#1 $display("%b", po);
# 1  pi=24'b010001101010001001111111;
#1 $display("%b", po);
# 1  pi=24'b100010101110001000100101;
#1 $display("%b", po);
# 1  pi=24'b000101100111000100000011;
#1 $display("%b", po);
# 1  pi=24'b000001101001010000100010;
#1 $display("%b", po);
# 1  pi=24'b000001000101111100101100;
#1 $display("%b", po);
# 1  pi=24'b110011010101100100101111;
#1 $display("%b", po);
# 1  pi=24'b001100010010000011001100;
#1 $display("%b", po);
# 1  pi=24'b111010001100011011111011;
#1 $display("%b", po);
# 1  pi=24'b011101011110010011101011;
#1 $display("%b", po);
# 1  pi=24'b100110110101110001111001;
#1 $display("%b", po);
# 1  pi=24'b100010111011010110110001;
#1 $display("%b", po);
# 1  pi=24'b011110111001011110010011;
#1 $display("%b", po);
# 1  pi=24'b010110110011001010001011;
#1 $display("%b", po);
# 1  pi=24'b111101100001001111101001;
#1 $display("%b", po);
# 1  pi=24'b001011100100000110100111;
#1 $display("%b", po);
# 1  pi=24'b111000011111110000000110;
#1 $display("%b", po);
# 1  pi=24'b010001001001101000011110;
#1 $display("%b", po);
# 1  pi=24'b111101101110100111101101;
#1 $display("%b", po);
# 1  pi=24'b111000001101110000100101;
#1 $display("%b", po);
# 1  pi=24'b101101001100000010010011;
#1 $display("%b", po);
# 1  pi=24'b100101101000110000100000;
#1 $display("%b", po);
# 1  pi=24'b111101110001011100011001;
#1 $display("%b", po);
# 1  pi=24'b111100011010010110001110;
#1 $display("%b", po);
# 1  pi=24'b101000010000000111100100;
#1 $display("%b", po);
# 1  pi=24'b000110111100010100110101;
#1 $display("%b", po);
# 1  pi=24'b110001101110100010100000;
#1 $display("%b", po);
# 1  pi=24'b011111111010000101111100;
#1 $display("%b", po);
# 1  pi=24'b010111011110111011111000;
#1 $display("%b", po);
# 1  pi=24'b101001010100111101110001;
#1 $display("%b", po);
# 1  pi=24'b110101011100001111000001;
#1 $display("%b", po);
# 1  pi=24'b100010011011010110001110;
#1 $display("%b", po);
# 1  pi=24'b001001011110101010000001;
#1 $display("%b", po);
# 1  pi=24'b111101011111010100101110;
#1 $display("%b", po);
# 1  pi=24'b011010100100011100000000;
#1 $display("%b", po);
# 1  pi=24'b001100100000001001100101;
#1 $display("%b", po);
# 1  pi=24'b000110110010100100001101;
#1 $display("%b", po);
# 1  pi=24'b000101011010100111110111;
#1 $display("%b", po);
# 1  pi=24'b010100001100111111011001;
#1 $display("%b", po);
# 1  pi=24'b000010110000111000111111;
#1 $display("%b", po);
# 1  pi=24'b000000101111001010101010;
#1 $display("%b", po);
# 1  pi=24'b101010111101011001000111;
#1 $display("%b", po);
# 1  pi=24'b011100011001011011101001;
#1 $display("%b", po);
# 1  pi=24'b101110110010001010010100;
#1 $display("%b", po);
# 1  pi=24'b011101011011010110111110;
#1 $display("%b", po);
# 1  pi=24'b100011000101000001001010;
#1 $display("%b", po);
# 1  pi=24'b101010010010111010010100;
#1 $display("%b", po);
# 1  pi=24'b110100110010101010011010;
#1 $display("%b", po);
# 1  pi=24'b001100010111111111100111;
#1 $display("%b", po);
# 1  pi=24'b100101011101010000101100;
#1 $display("%b", po);
# 1  pi=24'b011000001100100110100100;
#1 $display("%b", po);
# 1  pi=24'b101001110111111011110000;
#1 $display("%b", po);
# 1  pi=24'b001111110100111011100001;
#1 $display("%b", po);
# 1  pi=24'b001100011100111101001111;
#1 $display("%b", po);
# 1  pi=24'b000011110000011111101011;
#1 $display("%b", po);
# 1  pi=24'b111101110110001001101000;
#1 $display("%b", po);
# 1  pi=24'b010010010010111110101010;
#1 $display("%b", po);
# 1  pi=24'b001100011001110011010010;
#1 $display("%b", po);
# 1  pi=24'b100110001111010101110000;
#1 $display("%b", po);
# 1  pi=24'b001001111110100010101011;
#1 $display("%b", po);
# 1  pi=24'b111011100010101101111111;
#1 $display("%b", po);
# 1  pi=24'b000100100110100110011001;
#1 $display("%b", po);
# 1  pi=24'b110011011100010011001011;
#1 $display("%b", po);
# 1  pi=24'b001100111010011101100110;
#1 $display("%b", po);
# 1  pi=24'b100111000100100010010001;
#1 $display("%b", po);
# 1  pi=24'b101111011110111110010100;
#1 $display("%b", po);
# 1  pi=24'b011111000011101011100000;
#1 $display("%b", po);
# 1  pi=24'b111001101110101111111010;
#1 $display("%b", po);
# 1  pi=24'b001011011110111100101001;
#1 $display("%b", po);
# 1  pi=24'b101111011110000001101000;
#1 $display("%b", po);
# 1  pi=24'b101110110011000100001111;
#1 $display("%b", po);
# 1  pi=24'b001011101001000001001101;
#1 $display("%b", po);
# 1  pi=24'b000110011111011001000001;
#1 $display("%b", po);
# 1  pi=24'b100110000101100011010001;
#1 $display("%b", po);
# 1  pi=24'b110011001110001101011001;
#1 $display("%b", po);
# 1  pi=24'b101010111101010101000100;
#1 $display("%b", po);
# 1  pi=24'b110101101111010111111001;
#1 $display("%b", po);
# 1  pi=24'b100100000000011000010100;
#1 $display("%b", po);
# 1  pi=24'b011010110010010000010111;
#1 $display("%b", po);
# 1  pi=24'b101010110001110111100101;
#1 $display("%b", po);
# 1  pi=24'b101000111110011000100000;
#1 $display("%b", po);
# 1  pi=24'b001111100011100111001001;
#1 $display("%b", po);
# 1  pi=24'b001011110010001100110111;
#1 $display("%b", po);
# 1  pi=24'b011001111001110010111101;
#1 $display("%b", po);
# 1  pi=24'b011101001000011010000101;
#1 $display("%b", po);
# 1  pi=24'b001011110110010110010100;
#1 $display("%b", po);
# 1  pi=24'b001100110101111010000111;
#1 $display("%b", po);
# 1  pi=24'b010001010000000001010111;
#1 $display("%b", po);
# 1  pi=24'b000010100000100001101111;
#1 $display("%b", po);
# 1  pi=24'b001100011000001101001001;
#1 $display("%b", po);
# 1  pi=24'b011000010010001101001010;
#1 $display("%b", po);
# 1  pi=24'b111110010010001100101111;
#1 $display("%b", po);
# 1  pi=24'b000010000111101001011000;
#1 $display("%b", po);
# 1  pi=24'b101001000111100100000110;
#1 $display("%b", po);
# 1  pi=24'b001001000110111100010111;
#1 $display("%b", po);
# 1  pi=24'b000100101010011110110100;
#1 $display("%b", po);
# 1  pi=24'b110110000100001011001111;
#1 $display("%b", po);
# 1  pi=24'b010111100111000111110100;
#1 $display("%b", po);
# 1  pi=24'b010111101000011010110000;
#1 $display("%b", po);
# 1  pi=24'b001010111010100111001111;
#1 $display("%b", po);
# 1  pi=24'b110100010001111100101100;
#1 $display("%b", po);
# 1  pi=24'b111000001110111000000101;
#1 $display("%b", po);
# 1  pi=24'b000101000011100101010111;
#1 $display("%b", po);
# 1  pi=24'b000000110011000000011100;
#1 $display("%b", po);
# 1  pi=24'b101110101011100001001110;
#1 $display("%b", po);
# 1  pi=24'b111000010111110110110100;
#1 $display("%b", po);
# 1  pi=24'b010011001101101100111001;
#1 $display("%b", po);
# 1  pi=24'b000000111011011010010000;
#1 $display("%b", po);
# 1  pi=24'b001010010100000001000001;
#1 $display("%b", po);
# 1  pi=24'b110001010001010011111000;
#1 $display("%b", po);
# 1  pi=24'b110101111001011101001111;
#1 $display("%b", po);
# 1  pi=24'b111011011000101011001100;
#1 $display("%b", po);
# 1  pi=24'b110000001101001100000000;
#1 $display("%b", po);
# 1  pi=24'b111011010111101001010101;
#1 $display("%b", po);
# 1  pi=24'b110011010010101101101011;
#1 $display("%b", po);
# 1  pi=24'b111011100100010011011100;
#1 $display("%b", po);
# 1  pi=24'b110011010011001101010011;
#1 $display("%b", po);
# 1  pi=24'b010111101111110001010100;
#1 $display("%b", po);
# 1  pi=24'b100011010011111001000010;
#1 $display("%b", po);
# 1  pi=24'b111110100000000010011000;
#1 $display("%b", po);
# 1  pi=24'b000110110111100001001000;
#1 $display("%b", po);
# 1  pi=24'b100100111100001110100011;
#1 $display("%b", po);
# 1  pi=24'b100110100101001111100001;
#1 $display("%b", po);
# 1  pi=24'b011000110110100111010001;
#1 $display("%b", po);
# 1  pi=24'b010101010010010101110011;
#1 $display("%b", po);
# 1  pi=24'b101101010110100111000000;
#1 $display("%b", po);
# 1  pi=24'b100110101010100100111110;
#1 $display("%b", po);
# 1  pi=24'b110110111001000110000010;
#1 $display("%b", po);
# 1  pi=24'b101111001010100110001111;
#1 $display("%b", po);
# 1  pi=24'b100000010111000011010100;
#1 $display("%b", po);
# 1  pi=24'b011011010100000011111011;
#1 $display("%b", po);
# 1  pi=24'b111110110001110110110000;
#1 $display("%b", po);
# 1  pi=24'b101111110001110100011110;
#1 $display("%b", po);
# 1  pi=24'b110010001111011010010011;
#1 $display("%b", po);
# 1  pi=24'b001101001100110011000111;
#1 $display("%b", po);
# 1  pi=24'b100101001000010010100111;
#1 $display("%b", po);
# 1  pi=24'b110101101011111010101000;
#1 $display("%b", po);
# 1  pi=24'b100000100000001101110001;
#1 $display("%b", po);
# 1  pi=24'b101100110110011000100110;
#1 $display("%b", po);
# 1  pi=24'b011110010010010000010111;
#1 $display("%b", po);
# 1  pi=24'b111101110011010101011001;
#1 $display("%b", po);
# 1  pi=24'b010010011000010100101001;
#1 $display("%b", po);
# 1  pi=24'b111010011110101100010110;
#1 $display("%b", po);
# 1  pi=24'b000100000011001011101011;
#1 $display("%b", po);
# 1  pi=24'b000001011001001101000001;
#1 $display("%b", po);
# 1  pi=24'b001110000001101001110100;
#1 $display("%b", po);
# 1  pi=24'b001110110101001001010001;
#1 $display("%b", po);
# 1  pi=24'b010000011000101001001000;
#1 $display("%b", po);
# 1  pi=24'b000101111100111000011000;
#1 $display("%b", po);
# 1  pi=24'b010100010011100000111100;
#1 $display("%b", po);
# 1  pi=24'b110111100010001101100001;
#1 $display("%b", po);
# 1  pi=24'b111110101000101110000111;
#1 $display("%b", po);
# 1  pi=24'b101011110110110100110001;
#1 $display("%b", po);
# 1  pi=24'b000000001111000101011111;
#1 $display("%b", po);
# 1  pi=24'b011010100111010000100110;
#1 $display("%b", po);
# 1  pi=24'b101100111010100101111010;
#1 $display("%b", po);
# 1  pi=24'b011110111110001001010001;
#1 $display("%b", po);
# 1  pi=24'b110000101011010001010101;
#1 $display("%b", po);
# 1  pi=24'b110001001010110000011111;
#1 $display("%b", po);
# 1  pi=24'b001000101001000000101001;
#1 $display("%b", po);
# 1  pi=24'b101001111001111111111000;
#1 $display("%b", po);
# 1  pi=24'b101000001001100100011000;
#1 $display("%b", po);
# 1  pi=24'b100010111110000010001101;
#1 $display("%b", po);
# 1  pi=24'b110010010111011001100101;
#1 $display("%b", po);
# 1  pi=24'b111010001001000001011010;
#1 $display("%b", po);
# 1  pi=24'b111000110000110001110010;
#1 $display("%b", po);
# 1  pi=24'b110111001111110011111011;
#1 $display("%b", po);
# 1  pi=24'b000111101111011001111000;
#1 $display("%b", po);
# 1  pi=24'b001010000100011100110100;
#1 $display("%b", po);
# 1  pi=24'b011010111110011001110110;
#1 $display("%b", po);
# 1  pi=24'b010101010111000110101001;
#1 $display("%b", po);
# 1  pi=24'b100001001001000110000110;
#1 $display("%b", po);
# 1  pi=24'b110101110111100001111011;
#1 $display("%b", po);
# 1  pi=24'b110001101001100101001000;
#1 $display("%b", po);
# 1  pi=24'b000001001100011001010110;
#1 $display("%b", po);
# 1  pi=24'b011001011100011110011110;
#1 $display("%b", po);
# 1  pi=24'b100100001001110011100100;
#1 $display("%b", po);
# 1  pi=24'b011111111100100001111100;
#1 $display("%b", po);
# 1  pi=24'b000010111111011010100000;
#1 $display("%b", po);
# 1  pi=24'b011001000100101110110101;
#1 $display("%b", po);
# 1  pi=24'b101011111000001100101000;
#1 $display("%b", po);
# 1  pi=24'b010100011100111010111010;
#1 $display("%b", po);
# 1  pi=24'b111011100001100101111110;
#1 $display("%b", po);
# 1  pi=24'b001010010101001000100101;
#1 $display("%b", po);
# 1  pi=24'b011001100011001111001001;
#1 $display("%b", po);
# 1  pi=24'b010011000000111111101110;
#1 $display("%b", po);
# 1  pi=24'b010000000001101100000100;
#1 $display("%b", po);
# 1  pi=24'b110000011001110010001010;
#1 $display("%b", po);
# 1  pi=24'b000110101001001000100000;
#1 $display("%b", po);
# 1  pi=24'b000011010110101000101100;
#1 $display("%b", po);
# 1  pi=24'b011010001000001001111101;
#1 $display("%b", po);
# 1  pi=24'b010101101000000010000101;
#1 $display("%b", po);
# 1  pi=24'b101101011111110110101010;
#1 $display("%b", po);
# 1  pi=24'b111100011101010010000010;
#1 $display("%b", po);
# 1  pi=24'b110000011001011000100110;
#1 $display("%b", po);
# 1  pi=24'b101001000010100110011011;
#1 $display("%b", po);
# 1  pi=24'b011001100101100101001010;
#1 $display("%b", po);
# 1  pi=24'b010011100110100010100010;
#1 $display("%b", po);
# 1  pi=24'b100101011110001011100111;
#1 $display("%b", po);
# 1  pi=24'b000001101111101110001011;
#1 $display("%b", po);
# 1  pi=24'b010001000110111001010000;
#1 $display("%b", po);
# 1  pi=24'b011111110011111011111110;
#1 $display("%b", po);
# 1  pi=24'b100001001000111011010111;
#1 $display("%b", po);
# 1  pi=24'b000110010100011110000101;
#1 $display("%b", po);
# 1  pi=24'b111001110001101010000011;
#1 $display("%b", po);
# 1  pi=24'b111101101111010000111010;
#1 $display("%b", po);
# 1  pi=24'b000000111000001111000110;
#1 $display("%b", po);
# 1  pi=24'b001100111100001110111111;
#1 $display("%b", po);
# 1  pi=24'b010100001001000011011010;
#1 $display("%b", po);
# 1  pi=24'b010001011110110110111001;
#1 $display("%b", po);
# 1  pi=24'b110111011100110111001101;
#1 $display("%b", po);
# 1  pi=24'b001110001111000000100001;
#1 $display("%b", po);
# 1  pi=24'b000101111011010010110101;
#1 $display("%b", po);
# 1  pi=24'b010100101001011111010001;
#1 $display("%b", po);
# 1  pi=24'b010000111110010110111011;
#1 $display("%b", po);
# 1  pi=24'b000000011110110000100001;
#1 $display("%b", po);
# 1  pi=24'b001001100000110110101111;
#1 $display("%b", po);
# 1  pi=24'b010000011101110011101001;
#1 $display("%b", po);
# 1  pi=24'b011011000011110111100110;
#1 $display("%b", po);
# 1  pi=24'b010010100000010100001011;
#1 $display("%b", po);
# 1  pi=24'b001001110000100000100001;
#1 $display("%b", po);
# 1  pi=24'b111100100110101010011011;
#1 $display("%b", po);
# 1  pi=24'b110110011100010001010001;
#1 $display("%b", po);
# 1  pi=24'b011011101010100000000110;
#1 $display("%b", po);
# 1  pi=24'b000011001010000111111111;
#1 $display("%b", po);
# 1  pi=24'b111110010011111010000100;
#1 $display("%b", po);
# 1  pi=24'b111110001001000000001111;
#1 $display("%b", po);
# 1  pi=24'b100101000101010010001101;
#1 $display("%b", po);
# 1  pi=24'b100001011001100000000101;
#1 $display("%b", po);
# 1  pi=24'b101010001000001000100001;
#1 $display("%b", po);
# 1  pi=24'b100010101001111010111001;
#1 $display("%b", po);
# 1  pi=24'b111000101110001001110011;
#1 $display("%b", po);
# 1  pi=24'b011101101111001111001110;
#1 $display("%b", po);
# 1  pi=24'b001000110110110001110110;
#1 $display("%b", po);
# 1  pi=24'b001100011110001111100010;
#1 $display("%b", po);
# 1  pi=24'b100000100001011110100111;
#1 $display("%b", po);
# 1  pi=24'b110101011011100111100010;
#1 $display("%b", po);
# 1  pi=24'b101000001010100100010111;
#1 $display("%b", po);
# 1  pi=24'b011100111011111000110110;
#1 $display("%b", po);
# 1  pi=24'b011010111001000011110000;
#1 $display("%b", po);
# 1  pi=24'b010011111011001001100101;
#1 $display("%b", po);
# 1  pi=24'b001010000000010111101001;
#1 $display("%b", po);
# 1  pi=24'b110000101011100111101101;
#1 $display("%b", po);
# 1  pi=24'b101101001001100111011110;
#1 $display("%b", po);
# 1  pi=24'b110010100110110001011001;
#1 $display("%b", po);
# 1  pi=24'b000000000111011110010000;
#1 $display("%b", po);
# 1  pi=24'b111001010010101110110010;
#1 $display("%b", po);
# 1  pi=24'b111110011100111110110011;
#1 $display("%b", po);
# 1  pi=24'b101001011110101100101010;
#1 $display("%b", po);
# 1  pi=24'b100100011010010111000101;
#1 $display("%b", po);
# 1  pi=24'b110010111011110011011110;
#1 $display("%b", po);
# 1  pi=24'b001010011001010111110011;
#1 $display("%b", po);
# 1  pi=24'b111011111100100100100101;
#1 $display("%b", po);
# 1  pi=24'b101000011001011101010001;
#1 $display("%b", po);
# 1  pi=24'b011011100000100001010011;
#1 $display("%b", po);
# 1  pi=24'b110011010100111000101011;
#1 $display("%b", po);
# 1  pi=24'b011001000110001111100011;
#1 $display("%b", po);
# 1  pi=24'b010010110000011001110101;
#1 $display("%b", po);
# 1  pi=24'b111111011011100100101011;
#1 $display("%b", po);
# 1  pi=24'b101001001010000011011000;
#1 $display("%b", po);
# 1  pi=24'b100100011010100101001110;
#1 $display("%b", po);
# 1  pi=24'b111001100111100001111101;
#1 $display("%b", po);
# 1  pi=24'b001001001000000011000010;
#1 $display("%b", po);
# 1  pi=24'b101110111010011000110111;
#1 $display("%b", po);
# 1  pi=24'b100101100111011100100011;
#1 $display("%b", po);
# 1  pi=24'b110101011110000110110101;
#1 $display("%b", po);
# 1  pi=24'b000100111100110010110111;
#1 $display("%b", po);
# 1  pi=24'b100001001010010010011101;
#1 $display("%b", po);
# 1  pi=24'b001101110100000110101010;
#1 $display("%b", po);
# 1  pi=24'b101110000111011110110001;
#1 $display("%b", po);
# 1  pi=24'b000001001100000100011100;
#1 $display("%b", po);
# 1  pi=24'b101001010010110101110001;
#1 $display("%b", po);
# 1  pi=24'b101101011100011111100110;
#1 $display("%b", po);
# 1  pi=24'b011010110011011111101010;
#1 $display("%b", po);
# 1  pi=24'b101100111001100001001111;
#1 $display("%b", po);
# 1  pi=24'b101110010011110010000001;
#1 $display("%b", po);
# 1  pi=24'b000111101111001001110111;
#1 $display("%b", po);
# 1  pi=24'b010001110011010010111111;
#1 $display("%b", po);
# 1  pi=24'b001001011100010011110010;
#1 $display("%b", po);
# 1  pi=24'b010000111010011000101001;
#1 $display("%b", po);
# 1  pi=24'b011011001000001001111110;
#1 $display("%b", po);
# 1  pi=24'b100001000100000100011000;
#1 $display("%b", po);
# 1  pi=24'b000111000000101000011001;
#1 $display("%b", po);
# 1  pi=24'b101101010101111101010011;
#1 $display("%b", po);
# 1  pi=24'b010101101100111110000011;
#1 $display("%b", po);
# 1  pi=24'b111101100110010101000101;
#1 $display("%b", po);
# 1  pi=24'b011101111111010001110110;
#1 $display("%b", po);
# 1  pi=24'b101001110000100011100110;
#1 $display("%b", po);
# 1  pi=24'b111110001001100000001101;
#1 $display("%b", po);
# 1  pi=24'b101010101101110000100100;
#1 $display("%b", po);
# 1  pi=24'b101001101001111110111001;
#1 $display("%b", po);
# 1  pi=24'b000000101010010110100100;
#1 $display("%b", po);
# 1  pi=24'b100001111101011000100100;
#1 $display("%b", po);
# 1  pi=24'b010010011010011010100110;
#1 $display("%b", po);
# 1  pi=24'b101110111000101000011100;
#1 $display("%b", po);
# 1  pi=24'b001110101101001000010110;
#1 $display("%b", po);
# 1  pi=24'b001100000111111101001101;
#1 $display("%b", po);
# 1  pi=24'b010000111001111101110100;
#1 $display("%b", po);
# 1  pi=24'b101011101010010100100001;
#1 $display("%b", po);
# 1  pi=24'b001101100010100011101000;
#1 $display("%b", po);
# 1  pi=24'b010101110010110001010101;
#1 $display("%b", po);
# 1  pi=24'b010010000111000101101111;
#1 $display("%b", po);
# 1  pi=24'b000011001101001011011011;
#1 $display("%b", po);
# 1  pi=24'b011110010101000011010011;
#1 $display("%b", po);
# 1  pi=24'b001001111101001101110001;
#1 $display("%b", po);
# 1  pi=24'b111000001100110001101001;
#1 $display("%b", po);
# 1  pi=24'b101110100110011000101000;
#1 $display("%b", po);
# 1  pi=24'b111001111001000111010010;
#1 $display("%b", po);
# 1  pi=24'b110010110100010001000000;
#1 $display("%b", po);
# 1  pi=24'b100100101101011000100110;
#1 $display("%b", po);
# 1  pi=24'b100111111111100111101111;
#1 $display("%b", po);
# 1  pi=24'b110111100110011100101100;
#1 $display("%b", po);
# 1  pi=24'b001000001011110011010011;
#1 $display("%b", po);
# 1  pi=24'b110010111001110001110000;
#1 $display("%b", po);
# 1  pi=24'b000101000101001101010011;
#1 $display("%b", po);
# 1  pi=24'b110011110111101001000010;
#1 $display("%b", po);
# 1  pi=24'b001110001101001110111000;
#1 $display("%b", po);
# 1  pi=24'b011001011100100010011100;
#1 $display("%b", po);
# 1  pi=24'b101111111000011101001011;
#1 $display("%b", po);
# 1  pi=24'b001101111000010111101001;
#1 $display("%b", po);
# 1  pi=24'b101101110001000101110111;
#1 $display("%b", po);
# 1  pi=24'b101011101100101110101001;
#1 $display("%b", po);
# 1  pi=24'b111101111111100101000000;
#1 $display("%b", po);
# 1  pi=24'b011011001010111110001010;
#1 $display("%b", po);
# 1  pi=24'b100100101111010010010000;
#1 $display("%b", po);
# 1  pi=24'b100101100000111101001011;
#1 $display("%b", po);
# 1  pi=24'b000000001010100011001001;
#1 $display("%b", po);
# 1  pi=24'b001010010100111010111011;
#1 $display("%b", po);
# 1  pi=24'b100101100100000001010110;
#1 $display("%b", po);
# 1  pi=24'b001000001011100010101001;
#1 $display("%b", po);
# 1  pi=24'b100010111110101000101011;
#1 $display("%b", po);
# 1  pi=24'b011101010110011110011110;
#1 $display("%b", po);
# 1  pi=24'b011010010011010111011010;
#1 $display("%b", po);
# 1  pi=24'b000100111100101010110011;
#1 $display("%b", po);
# 1  pi=24'b011111011010000011111110;
#1 $display("%b", po);
# 1  pi=24'b000001100000101011101001;
#1 $display("%b", po);
# 1  pi=24'b100111001111101111101101;
#1 $display("%b", po);
# 1  pi=24'b110011000011101101011100;
#1 $display("%b", po);
# 1  pi=24'b000110000100000001010010;
#1 $display("%b", po);
# 1  pi=24'b101001100110110101010011;
#1 $display("%b", po);
# 1  pi=24'b000111000001010110001000;
#1 $display("%b", po);
# 1  pi=24'b011111100111000101011100;
#1 $display("%b", po);
# 1  pi=24'b110010110111011010001101;
#1 $display("%b", po);
# 1  pi=24'b011100000111000010001000;
#1 $display("%b", po);
# 1  pi=24'b011010111011000100110010;
#1 $display("%b", po);
# 1  pi=24'b000110111100110011100011;
#1 $display("%b", po);
# 1  pi=24'b110101100010001111011010;
#1 $display("%b", po);
# 1  pi=24'b100101110010100010010000;
#1 $display("%b", po);
# 1  pi=24'b110000001001000001111111;
#1 $display("%b", po);
# 1  pi=24'b100001001001100111101110;
#1 $display("%b", po);
# 1  pi=24'b111110110001001010111010;
#1 $display("%b", po);
# 1  pi=24'b101101111011000100001010;
#1 $display("%b", po);
# 1  pi=24'b010111110010010101010011;
#1 $display("%b", po);
# 1  pi=24'b110000110111001101000100;
#1 $display("%b", po);
# 1  pi=24'b111001100110001000100100;
#1 $display("%b", po);
# 1  pi=24'b001001110000101000101111;
#1 $display("%b", po);
# 1  pi=24'b100001010100101110111010;
#1 $display("%b", po);
# 1  pi=24'b110110010001001000111001;
#1 $display("%b", po);
# 1  pi=24'b001011101100011110010001;
#1 $display("%b", po);
# 1  pi=24'b110010111001001000011001;
#1 $display("%b", po);
# 1  pi=24'b110011010111110000000000;
#1 $display("%b", po);
# 1  pi=24'b011110111001000111000100;
#1 $display("%b", po);
# 1  pi=24'b001100110000001001011010;
#1 $display("%b", po);
# 1  pi=24'b111001000111111111100011;
#1 $display("%b", po);
# 1  pi=24'b100010001111110110100111;
#1 $display("%b", po);
# 1  pi=24'b111111010010100111110010;
#1 $display("%b", po);
# 1  pi=24'b010111011111010010010100;
#1 $display("%b", po);
# 1  pi=24'b011000111111011111001010;
#1 $display("%b", po);
# 1  pi=24'b111000111111011010110010;
#1 $display("%b", po);
# 1  pi=24'b100001000100011100010101;
#1 $display("%b", po);
# 1  pi=24'b100011001010100000011101;
#1 $display("%b", po);
# 1  pi=24'b100001011110111000000110;
#1 $display("%b", po);
# 1  pi=24'b011011011100000111010010;
#1 $display("%b", po);
# 1  pi=24'b100010001100101100110001;
#1 $display("%b", po);
# 1  pi=24'b011010000110111010001001;
#1 $display("%b", po);
# 1  pi=24'b101111011100111110101010;
#1 $display("%b", po);
# 1  pi=24'b100011100000110010100001;
#1 $display("%b", po);
# 1  pi=24'b100100111110110001000001;
#1 $display("%b", po);
# 1  pi=24'b110100010001111011111101;
#1 $display("%b", po);
# 1  pi=24'b111111000000011000011011;
#1 $display("%b", po);
# 1  pi=24'b011010110010001001011110;
#1 $display("%b", po);
# 1  pi=24'b010001110010000001000111;
#1 $display("%b", po);
# 1  pi=24'b001110001110011001100001;
#1 $display("%b", po);
# 1  pi=24'b101101010000100101100011;
#1 $display("%b", po);
# 1  pi=24'b111001000100101011001000;
#1 $display("%b", po);
# 1  pi=24'b010010010011001000100000;
#1 $display("%b", po);
# 1  pi=24'b100101100000110100111111;
#1 $display("%b", po);
# 1  pi=24'b000100101101010010110000;
#1 $display("%b", po);
# 1  pi=24'b011001101110110010101001;
#1 $display("%b", po);
# 1  pi=24'b011011001110011010100111;
#1 $display("%b", po);
# 1  pi=24'b001111110110100001101111;
#1 $display("%b", po);
# 1  pi=24'b000111111000100110101011;
#1 $display("%b", po);
# 1  pi=24'b011001000011110011010101;
#1 $display("%b", po);
# 1  pi=24'b111110010001010110011111;
#1 $display("%b", po);
# 1  pi=24'b000000100100010101100001;
#1 $display("%b", po);
# 1  pi=24'b001100001110111010011000;
#1 $display("%b", po);
# 1  pi=24'b001010101100110001010110;
#1 $display("%b", po);
# 1  pi=24'b111100010101010000010100;
#1 $display("%b", po);
# 1  pi=24'b110001000100100100101011;
#1 $display("%b", po);
# 1  pi=24'b100110000110111010111011;
#1 $display("%b", po);
# 1  pi=24'b010101111100111110101100;
#1 $display("%b", po);
# 1  pi=24'b010100100010010111111111;
#1 $display("%b", po);
# 1  pi=24'b010010101011001010001000;
#1 $display("%b", po);
# 1  pi=24'b110101101011010100000110;
#1 $display("%b", po);
# 1  pi=24'b001000010111101010001110;
#1 $display("%b", po);
# 1  pi=24'b111101111000101011100001;
#1 $display("%b", po);
# 1  pi=24'b110111101000110111100100;
#1 $display("%b", po);
# 1  pi=24'b010101001000111000001010;
#1 $display("%b", po);
# 1  pi=24'b011010001001100110010010;
#1 $display("%b", po);
# 1  pi=24'b000010111101000000010110;
#1 $display("%b", po);
# 1  pi=24'b101100011100011011110000;
#1 $display("%b", po);
# 1  pi=24'b100001001110000110001000;
#1 $display("%b", po);
# 1  pi=24'b111000000101000011010011;
#1 $display("%b", po);
# 1  pi=24'b100111111001010100011110;
#1 $display("%b", po);
# 1  pi=24'b001010111001001101110000;
#1 $display("%b", po);
# 1  pi=24'b011011111110100111000110;
#1 $display("%b", po);
# 1  pi=24'b000101100011000001010000;
#1 $display("%b", po);
# 1  pi=24'b000010111100111011100010;
#1 $display("%b", po);
# 1  pi=24'b010100000000101010101111;
#1 $display("%b", po);
# 1  pi=24'b010110000111011011111111;
#1 $display("%b", po);
# 1  pi=24'b110010100101100111101111;
#1 $display("%b", po);
# 1  pi=24'b011010011011011111001111;
#1 $display("%b", po);
# 1  pi=24'b100010111000011011100111;
#1 $display("%b", po);
# 1  pi=24'b000011110000011110110000;
#1 $display("%b", po);
# 1  pi=24'b001001000000000111100111;
#1 $display("%b", po);
# 1  pi=24'b010110100001101110111011;
#1 $display("%b", po);
# 1  pi=24'b001101000100010001001011;
#1 $display("%b", po);
# 1  pi=24'b110001110011011111110010;
#1 $display("%b", po);
# 1  pi=24'b111010100011011000000000;
#1 $display("%b", po);
# 1  pi=24'b001110101010101001011010;
#1 $display("%b", po);
# 1  pi=24'b101001010111001101110100;
#1 $display("%b", po);
# 1  pi=24'b001111000000010011101010;
#1 $display("%b", po);
# 1  pi=24'b010000100110110011100100;
#1 $display("%b", po);
# 1  pi=24'b010001010111000001010100;
#1 $display("%b", po);
# 1  pi=24'b100100000101011011110011;
#1 $display("%b", po);
# 1  pi=24'b001101111100110001101001;
#1 $display("%b", po);
# 1  pi=24'b100000001011001000011010;
#1 $display("%b", po);
# 1  pi=24'b010010101001010010100000;
#1 $display("%b", po);
# 1  pi=24'b111101111010010110111010;
#1 $display("%b", po);
# 1  pi=24'b110001010010001010000011;
#1 $display("%b", po);
# 1  pi=24'b110111001100001101000000;
#1 $display("%b", po);
# 1  pi=24'b011010100001011011000100;
#1 $display("%b", po);
# 1  pi=24'b000101101000001101000100;
#1 $display("%b", po);
# 1  pi=24'b111111001110110000100101;
#1 $display("%b", po);
# 1  pi=24'b010000101001000110011010;
#1 $display("%b", po);
# 1  pi=24'b010111101000001010011101;
#1 $display("%b", po);
# 1  pi=24'b000111001011100001111000;
#1 $display("%b", po);
# 1  pi=24'b001000100010011011101111;
#1 $display("%b", po);
# 1  pi=24'b000011101010000010111110;
#1 $display("%b", po);
# 1  pi=24'b000101110100010111000000;
#1 $display("%b", po);
# 1  pi=24'b000010110111000100000010;
#1 $display("%b", po);
# 1  pi=24'b011000011111101111101011;
#1 $display("%b", po);
# 1  pi=24'b101010110110111010011001;
#1 $display("%b", po);
# 1  pi=24'b001010001110010111111100;
#1 $display("%b", po);
# 1  pi=24'b110000101001101110111001;
#1 $display("%b", po);
# 1  pi=24'b110101000001000111101110;
#1 $display("%b", po);
# 1  pi=24'b011100010101111110100101;
#1 $display("%b", po);
# 1  pi=24'b000011000000110110101100;
#1 $display("%b", po);
# 1  pi=24'b010011100101011010111110;
#1 $display("%b", po);
# 1  pi=24'b110000100110000110011001;
#1 $display("%b", po);
# 1  pi=24'b011100010011111101100100;
#1 $display("%b", po);
# 1  pi=24'b110000100000011100011000;
#1 $display("%b", po);
# 1  pi=24'b100100011001110111100010;
#1 $display("%b", po);
# 1  pi=24'b111111011000001011100011;
#1 $display("%b", po);
# 1  pi=24'b001000100000110011100001;
#1 $display("%b", po);
# 1  pi=24'b011001101000110011011001;
#1 $display("%b", po);
# 1  pi=24'b111101100001101010111000;
#1 $display("%b", po);
# 1  pi=24'b101100011101101000000011;
#1 $display("%b", po);
# 1  pi=24'b110101000010010010100001;
#1 $display("%b", po);
# 1  pi=24'b110001001111001011110101;
#1 $display("%b", po);
# 1  pi=24'b010011100111111001011001;
#1 $display("%b", po);
# 1  pi=24'b000011101100000010010110;
#1 $display("%b", po);
# 1  pi=24'b110011011111110101100000;
#1 $display("%b", po);
# 1  pi=24'b001100000101011101010001;
#1 $display("%b", po);
# 1  pi=24'b100000010111101011000010;
#1 $display("%b", po);
# 1  pi=24'b001001010101111100101000;
#1 $display("%b", po);
# 1  pi=24'b000111111101101110101001;
#1 $display("%b", po);
# 1  pi=24'b010001110000000010110101;
#1 $display("%b", po);
# 1  pi=24'b001001011001000011100101;
#1 $display("%b", po);
# 1  pi=24'b000011111000110001100100;
#1 $display("%b", po);
# 1  pi=24'b111011000010001111010001;
#1 $display("%b", po);
# 1  pi=24'b101100100110101110101001;
#1 $display("%b", po);
# 1  pi=24'b001101010110010000110101;
#1 $display("%b", po);
# 1  pi=24'b000101110010110010000011;
#1 $display("%b", po);
# 1  pi=24'b101111011100101000000011;
#1 $display("%b", po);
# 1  pi=24'b010000000010010011011100;
#1 $display("%b", po);
# 1  pi=24'b001101000001001101101010;
#1 $display("%b", po);
# 1  pi=24'b110111000101001111100111;
#1 $display("%b", po);
# 1  pi=24'b111010101101010100101111;
#1 $display("%b", po);
# 1  pi=24'b100110001010011100101110;
#1 $display("%b", po);
# 1  pi=24'b111001110001101001100111;
#1 $display("%b", po);
# 1  pi=24'b101101101110001100001100;
#1 $display("%b", po);
# 1  pi=24'b111011100111111100010001;
#1 $display("%b", po);
# 1  pi=24'b111101100111101100110010;
#1 $display("%b", po);
# 1  pi=24'b000111001001111101111011;
#1 $display("%b", po);
# 1  pi=24'b100010110010111000010101;
#1 $display("%b", po);
# 1  pi=24'b011000000100111101010100;
#1 $display("%b", po);
# 1  pi=24'b011100001110110110000100;
#1 $display("%b", po);
# 1  pi=24'b101100010001111011001111;
#1 $display("%b", po);
# 1  pi=24'b010001110010010001010100;
#1 $display("%b", po);
# 1  pi=24'b010011000111000001111101;
#1 $display("%b", po);
# 1  pi=24'b100100101001100111011010;
#1 $display("%b", po);
# 1  pi=24'b110010000011110101010011;
#1 $display("%b", po);
# 1  pi=24'b011101101110110101110100;
#1 $display("%b", po);
# 1  pi=24'b100011100111111001010001;
#1 $display("%b", po);
# 1  pi=24'b101001010000011000100001;
#1 $display("%b", po);
# 1  pi=24'b100100101011011000011111;
#1 $display("%b", po);
# 1  pi=24'b010101011111011101011100;
#1 $display("%b", po);
# 1  pi=24'b011011101010100111001001;
#1 $display("%b", po);
# 1  pi=24'b000001100101111000010001;
#1 $display("%b", po);
# 1  pi=24'b101010010001100110101001;
#1 $display("%b", po);
# 1  pi=24'b111101111111101000010101;
#1 $display("%b", po);
# 1  pi=24'b000111111100011101110100;
#1 $display("%b", po);
# 1  pi=24'b000011011111100110010010;
#1 $display("%b", po);
# 1  pi=24'b010011110110110100100001;
#1 $display("%b", po);
# 1  pi=24'b011100000110000001001111;
#1 $display("%b", po);
# 1  pi=24'b100110101100100010110001;
#1 $display("%b", po);
# 1  pi=24'b000001100001100100101110;
#1 $display("%b", po);
# 1  pi=24'b100001010110010010010000;
#1 $display("%b", po);
# 1  pi=24'b111001111111111010011011;
#1 $display("%b", po);
# 1  pi=24'b100001010110110011001011;
#1 $display("%b", po);
# 1  pi=24'b011010010001100111000101;
#1 $display("%b", po);
# 1  pi=24'b101100011010000101001010;
#1 $display("%b", po);
# 1  pi=24'b001010111101001001111111;
#1 $display("%b", po);
# 1  pi=24'b111001110100000100010000;
#1 $display("%b", po);
# 1  pi=24'b011100011111010010010011;
#1 $display("%b", po);
# 1  pi=24'b100100110100011000100010;
#1 $display("%b", po);
# 1  pi=24'b100000000001011110111101;
#1 $display("%b", po);
# 1  pi=24'b110010110100100100000100;
#1 $display("%b", po);
# 1  pi=24'b010011110100001011001000;
#1 $display("%b", po);
# 1  pi=24'b110111100010110001011011;
#1 $display("%b", po);
# 1  pi=24'b101110111010010001111010;
#1 $display("%b", po);
# 1  pi=24'b001100110101101010110111;
#1 $display("%b", po);
# 1  pi=24'b101111110011001111001000;
#1 $display("%b", po);
# 1  pi=24'b001100000111000100001010;
#1 $display("%b", po);
# 1  pi=24'b001101100111101101101000;
#1 $display("%b", po);
# 1  pi=24'b111111000011000011100001;
#1 $display("%b", po);
# 1  pi=24'b000010101100000001100011;
#1 $display("%b", po);
# 1  pi=24'b100100001101110001010001;
#1 $display("%b", po);
# 1  pi=24'b111100000010111100010011;
#1 $display("%b", po);
# 1  pi=24'b001111001000001011111110;
#1 $display("%b", po);
# 1  pi=24'b111000101110001110111100;
#1 $display("%b", po);
# 1  pi=24'b100111001101001100101111;
#1 $display("%b", po);
# 1  pi=24'b111110101101100010101101;
#1 $display("%b", po);
# 1  pi=24'b000100100010110101101001;
#1 $display("%b", po);
# 1  pi=24'b010011100010000000001011;
#1 $display("%b", po);
# 1  pi=24'b000011111101000011011000;
#1 $display("%b", po);
# 1  pi=24'b011100000110101001000100;
#1 $display("%b", po);
# 1  pi=24'b100001100000101001101001;
#1 $display("%b", po);
# 1  pi=24'b011101110001001001000101;
#1 $display("%b", po);
# 1  pi=24'b111101110110100010001001;
#1 $display("%b", po);
# 1  pi=24'b010000110000100110110101;
#1 $display("%b", po);
# 1  pi=24'b110010011000100100101101;
#1 $display("%b", po);
# 1  pi=24'b010110101100010011101011;
#1 $display("%b", po);
# 1  pi=24'b011101100011001000100010;
#1 $display("%b", po);
# 1  pi=24'b110010111010011110001101;
#1 $display("%b", po);
# 1  pi=24'b010011110011101111110111;
#1 $display("%b", po);
# 1  pi=24'b111101000011001100100111;
#1 $display("%b", po);
# 1  pi=24'b001000000000111000010011;
#1 $display("%b", po);
# 1  pi=24'b100111000011101000100110;
#1 $display("%b", po);
# 1  pi=24'b100101111100100101011011;
#1 $display("%b", po);
# 1  pi=24'b001010001110011100000001;
#1 $display("%b", po);
# 1  pi=24'b010010110111011000111101;
#1 $display("%b", po);
# 1  pi=24'b100101110000001011010111;
#1 $display("%b", po);
# 1  pi=24'b011110111001001100100111;
#1 $display("%b", po);
# 1  pi=24'b100001010110000000001010;
#1 $display("%b", po);
# 1  pi=24'b111101011001100100111110;
#1 $display("%b", po);
# 1  pi=24'b110000101101001101000101;
#1 $display("%b", po);
# 1  pi=24'b001100111001101111000011;
#1 $display("%b", po);
# 1  pi=24'b111110011010110000010001;
#1 $display("%b", po);
# 1  pi=24'b000001100011011010100011;
#1 $display("%b", po);
# 1  pi=24'b101110110011101111011000;
#1 $display("%b", po);
# 1  pi=24'b000001111111001111010001;
#1 $display("%b", po);
# 1  pi=24'b010111111010101111100001;
#1 $display("%b", po);
# 1  pi=24'b110111000010100010001001;
#1 $display("%b", po);
# 1  pi=24'b100100100101010111000000;
#1 $display("%b", po);
# 1  pi=24'b011111110111001101101100;
#1 $display("%b", po);
# 1  pi=24'b111110101011111000011000;
#1 $display("%b", po);
# 1  pi=24'b000010101011001010100010;
#1 $display("%b", po);
# 1  pi=24'b111010101010101011010011;
#1 $display("%b", po);
# 1  pi=24'b100110001001111000000110;
#1 $display("%b", po);
# 1  pi=24'b001000010011101010000000;
#1 $display("%b", po);
# 1  pi=24'b101011011100011111001011;
#1 $display("%b", po);
# 1  pi=24'b010101111000101100101001;
#1 $display("%b", po);
# 1  pi=24'b011011111010110110000110;
#1 $display("%b", po);
# 1  pi=24'b100001101011011110100010;
#1 $display("%b", po);
# 1  pi=24'b010000111100000110011010;
#1 $display("%b", po);
# 1  pi=24'b010110111000110011101110;
#1 $display("%b", po);
# 1  pi=24'b100100101011001100010000;
#1 $display("%b", po);
# 1  pi=24'b101110111110001001101111;
#1 $display("%b", po);
# 1  pi=24'b111111001011101111110110;
#1 $display("%b", po);
# 1  pi=24'b110101010111000000101010;
#1 $display("%b", po);
# 1  pi=24'b011111011000000101000011;
#1 $display("%b", po);
# 1  pi=24'b101001110100001000010110;
#1 $display("%b", po);
# 1  pi=24'b011000000011110111101111;
#1 $display("%b", po);
# 1  pi=24'b010000101111000101110001;
#1 $display("%b", po);
# 1  pi=24'b000000001100111111100110;
#1 $display("%b", po);
# 1  pi=24'b110100111111111000101001;
#1 $display("%b", po);
# 1  pi=24'b010111010111100000010000;
#1 $display("%b", po);
# 1  pi=24'b010101110110100111101111;
#1 $display("%b", po);
# 1  pi=24'b000100111001001001101111;
#1 $display("%b", po);
# 1  pi=24'b100011000010000001111001;
#1 $display("%b", po);
# 1  pi=24'b010000100010100001011101;
#1 $display("%b", po);
# 1  pi=24'b000001000100000010000001;
#1 $display("%b", po);
# 1  pi=24'b000111110011111101100001;
#1 $display("%b", po);
# 1  pi=24'b100111010101101011111110;
#1 $display("%b", po);
# 1  pi=24'b011001100011101110011101;
#1 $display("%b", po);
# 1  pi=24'b110111000111011000011000;
#1 $display("%b", po);
# 1  pi=24'b101111110001010101101100;
#1 $display("%b", po);
# 1  pi=24'b011100011010110101110110;
#1 $display("%b", po);
# 1  pi=24'b010001001001001001000011;
#1 $display("%b", po);
# 1  pi=24'b000111111100001110011000;
#1 $display("%b", po);
# 1  pi=24'b111001111101100101101100;
#1 $display("%b", po);
# 1  pi=24'b101000101000011001101000;
#1 $display("%b", po);
# 1  pi=24'b010001001111101110010001;
#1 $display("%b", po);
# 1  pi=24'b110101010110000001110111;
#1 $display("%b", po);
# 1  pi=24'b011010101010001001111101;
#1 $display("%b", po);
# 1  pi=24'b000101001110111001010011;
#1 $display("%b", po);
# 1  pi=24'b101010110000001101101011;
#1 $display("%b", po);
# 1  pi=24'b010111001010010110111100;
#1 $display("%b", po);
# 1  pi=24'b100010000000001000001110;
#1 $display("%b", po);
# 1  pi=24'b110111001001011010111011;
#1 $display("%b", po);
# 1  pi=24'b010011100011011011011110;
#1 $display("%b", po);
# 1  pi=24'b111100110011011001010000;
#1 $display("%b", po);
# 1  pi=24'b011110110001011000000011;
#1 $display("%b", po);
# 1  pi=24'b000010110100001111101010;
#1 $display("%b", po);
# 1  pi=24'b011100111110111111010001;
#1 $display("%b", po);
# 1  pi=24'b000110000000001111011101;
#1 $display("%b", po);
# 1  pi=24'b011011110101110100000101;
#1 $display("%b", po);
# 1  pi=24'b001000100111001010111110;
#1 $display("%b", po);
# 1  pi=24'b000111011011100010011111;
#1 $display("%b", po);
# 1  pi=24'b011110011110110111111010;
#1 $display("%b", po);
# 1  pi=24'b010111000011000001110010;
#1 $display("%b", po);
# 1  pi=24'b011111100110010010010000;
#1 $display("%b", po);
# 1  pi=24'b011110101101110111100100;
#1 $display("%b", po);
# 1  pi=24'b010111111010001100101010;
#1 $display("%b", po);
# 1  pi=24'b000111011110000101110101;
#1 $display("%b", po);
# 1  pi=24'b000000000010001011000011;
#1 $display("%b", po);
# 1  pi=24'b110110011000110001110010;
#1 $display("%b", po);
# 1  pi=24'b000101110110001110011101;
#1 $display("%b", po);
# 1  pi=24'b010000100110001010100100;
#1 $display("%b", po);
# 1  pi=24'b111110011110101100111010;
#1 $display("%b", po);
# 1  pi=24'b000010001100001000011000;
#1 $display("%b", po);
# 1  pi=24'b011110100000001001111100;
#1 $display("%b", po);
# 1  pi=24'b010100000010011010000111;
#1 $display("%b", po);
# 1  pi=24'b001100111101111100001111;
#1 $display("%b", po);
# 1  pi=24'b110100001001011001110000;
#1 $display("%b", po);
# 1  pi=24'b001001101111110110011100;
#1 $display("%b", po);
# 1  pi=24'b011011100000111011001000;
#1 $display("%b", po);
# 1  pi=24'b101011000101111000001111;
#1 $display("%b", po);
# 1  pi=24'b101001100110011010101101;
#1 $display("%b", po);
# 1  pi=24'b001100100100101001111111;
#1 $display("%b", po);
# 1  pi=24'b101000100110100101000110;
#1 $display("%b", po);
# 1  pi=24'b111111010101110111101000;
#1 $display("%b", po);
# 1  pi=24'b000011000010101100010011;
#1 $display("%b", po);
# 1  pi=24'b100111000111000100100101;
#1 $display("%b", po);
# 1  pi=24'b111111111000001000100001;
#1 $display("%b", po);
# 1  pi=24'b110111110010000011110101;
#1 $display("%b", po);
# 1  pi=24'b010011100011000011111110;
#1 $display("%b", po);
# 1  pi=24'b110000000100100000001010;
#1 $display("%b", po);
# 1  pi=24'b101011100111011100101111;
#1 $display("%b", po);
# 1  pi=24'b010001011110001100001011;
#1 $display("%b", po);
# 1  pi=24'b111100010111000010010111;
#1 $display("%b", po);
# 1  pi=24'b111110011111101110011000;
#1 $display("%b", po);
# 1  pi=24'b000100000111000110101110;
#1 $display("%b", po);
# 1  pi=24'b010000111111110001111001;
#1 $display("%b", po);
# 1  pi=24'b000101011100100011110111;
#1 $display("%b", po);
# 1  pi=24'b101011111110000101011001;
#1 $display("%b", po);
# 1  pi=24'b011011101001010101010100;
#1 $display("%b", po);
# 1  pi=24'b110010001111001011000101;
#1 $display("%b", po);
# 1  pi=24'b011001101011000111101011;
#1 $display("%b", po);
# 1  pi=24'b110100111101001110111110;
#1 $display("%b", po);
# 1  pi=24'b000100101010101111001001;
#1 $display("%b", po);
# 1  pi=24'b001111011101001011101111;
#1 $display("%b", po);
# 1  pi=24'b010110101000000101011100;
#1 $display("%b", po);
# 1  pi=24'b001111101011001101000001;
#1 $display("%b", po);
# 1  pi=24'b110101110001100101011010;
#1 $display("%b", po);
# 1  pi=24'b010001000010001110010000;
#1 $display("%b", po);
# 1  pi=24'b011000111001110010000111;
#1 $display("%b", po);
# 1  pi=24'b010001110101111010111110;
#1 $display("%b", po);
# 1  pi=24'b011111011010101110110010;
#1 $display("%b", po);
# 1  pi=24'b010010100111110111100111;
#1 $display("%b", po);
# 1  pi=24'b010101100011001110100000;
#1 $display("%b", po);
# 1  pi=24'b011001111010000101100010;
#1 $display("%b", po);
# 1  pi=24'b111111101011010110111000;
#1 $display("%b", po);
# 1  pi=24'b101101111011010100000101;
#1 $display("%b", po);
# 1  pi=24'b010010100001100110110010;
#1 $display("%b", po);
# 1  pi=24'b000101101000001110100101;
#1 $display("%b", po);
# 1  pi=24'b001100100100111000111101;
#1 $display("%b", po);
# 1  pi=24'b111110011011110011101101;
#1 $display("%b", po);
# 1  pi=24'b001011000111001010111100;
#1 $display("%b", po);
# 1  pi=24'b010000101011111111001000;
#1 $display("%b", po);
# 1  pi=24'b010101010101110000010001;
#1 $display("%b", po);
# 1  pi=24'b101011010100111101111110;
#1 $display("%b", po);
# 1  pi=24'b110000100010000011111101;
#1 $display("%b", po);
# 1  pi=24'b000100100011000111111110;
#1 $display("%b", po);
# 1  pi=24'b000000001010010000111110;
#1 $display("%b", po);
# 1  pi=24'b101001110111111110111101;
#1 $display("%b", po);
# 1  pi=24'b110111111101010001111001;
#1 $display("%b", po);
# 1  pi=24'b001001111010010111000000;
#1 $display("%b", po);
# 1  pi=24'b001100100010100011101111;
#1 $display("%b", po);
# 1  pi=24'b011101111011000001000000;
#1 $display("%b", po);
# 1  pi=24'b000000110100111001010111;
#1 $display("%b", po);
# 1  pi=24'b011000101100011101001111;
#1 $display("%b", po);
# 1  pi=24'b100001110100011001100101;
#1 $display("%b", po);
# 1  pi=24'b101001100101110101111101;
#1 $display("%b", po);
# 1  pi=24'b110100110001010101011101;
#1 $display("%b", po);
# 1  pi=24'b100110100110111000100111;
#1 $display("%b", po);
# 1  pi=24'b100011110110111010100010;
#1 $display("%b", po);
# 1  pi=24'b101100010100000001001110;
#1 $display("%b", po);
# 1  pi=24'b110011111111111010000111;
#1 $display("%b", po);
# 1  pi=24'b101010000011011010001110;
#1 $display("%b", po);
# 1  pi=24'b101010101110010011110001;
#1 $display("%b", po);
# 1  pi=24'b001111100111111110110111;
#1 $display("%b", po);
# 1  pi=24'b011100011010110101110000;
#1 $display("%b", po);
# 1  pi=24'b101011111011000101111010;
#1 $display("%b", po);
# 1  pi=24'b101101111111011111001110;
#1 $display("%b", po);
# 1  pi=24'b100010001110001011111111;
#1 $display("%b", po);
# 1  pi=24'b110110111110000101011111;
#1 $display("%b", po);
# 1  pi=24'b101110111100011100101001;
#1 $display("%b", po);
# 1  pi=24'b010000111011010101010001;
#1 $display("%b", po);
# 1  pi=24'b011110100100000110001000;
#1 $display("%b", po);
# 1  pi=24'b010000111101011001000001;
#1 $display("%b", po);
# 1  pi=24'b101110100111000010101010;
#1 $display("%b", po);
# 1  pi=24'b001000100110011010110101;
#1 $display("%b", po);
# 1  pi=24'b010001110000011111101111;
#1 $display("%b", po);
# 1  pi=24'b000101001010110110110101;
#1 $display("%b", po);
# 1  pi=24'b100010000011100100110001;
#1 $display("%b", po);
# 1  pi=24'b110000100011110101110000;
#1 $display("%b", po);
# 1  pi=24'b010010100000111110011000;
#1 $display("%b", po);
# 1  pi=24'b000011000111001101101001;
#1 $display("%b", po);
# 1  pi=24'b101011000001110111000001;
#1 $display("%b", po);
# 1  pi=24'b111101001010100010001100;
#1 $display("%b", po);
# 1  pi=24'b011001001000001010111000;
#1 $display("%b", po);
# 1  pi=24'b010101100111011111100101;
#1 $display("%b", po);
# 1  pi=24'b001000000111011001100010;
#1 $display("%b", po);
# 1  pi=24'b111001110011110011100111;
#1 $display("%b", po);
# 1  pi=24'b100010101010011110111011;
#1 $display("%b", po);
# 1  pi=24'b110110011100011110100111;
#1 $display("%b", po);
# 1  pi=24'b111111010010110110010000;
#1 $display("%b", po);
# 1  pi=24'b000100010100011010011100;
#1 $display("%b", po);
# 1  pi=24'b011010101101101011000111;
#1 $display("%b", po);
# 1  pi=24'b111010110110101111100010;
#1 $display("%b", po);
# 1  pi=24'b110111000100001001000110;
#1 $display("%b", po);
# 1  pi=24'b010100110101100111011011;
#1 $display("%b", po);
# 1  pi=24'b010111111010111100011000;
#1 $display("%b", po);
# 1  pi=24'b100010101000100010010101;
#1 $display("%b", po);
# 1  pi=24'b011111100100001111010010;
#1 $display("%b", po);
# 1  pi=24'b110011100100111000001001;
#1 $display("%b", po);
# 1  pi=24'b010011110100110010101110;
#1 $display("%b", po);
# 1  pi=24'b111000111011101000111010;
#1 $display("%b", po);
# 1  pi=24'b011100010111011011001010;
#1 $display("%b", po);
# 1  pi=24'b000111111001111001001010;
#1 $display("%b", po);
# 1  pi=24'b110010110000010110111011;
#1 $display("%b", po);
# 1  pi=24'b110011001000101111011001;
#1 $display("%b", po);
# 1  pi=24'b010001000000001001001011;
#1 $display("%b", po);
# 1  pi=24'b101011011101111001000111;
#1 $display("%b", po);
# 1  pi=24'b111101001001010110001111;
#1 $display("%b", po);
# 1  pi=24'b011011110111110111011011;
#1 $display("%b", po);
# 1  pi=24'b010101101100101100010100;
#1 $display("%b", po);
# 1  pi=24'b111011000011000100110011;
#1 $display("%b", po);
# 1  pi=24'b010110111000110010100000;
#1 $display("%b", po);
# 1  pi=24'b000001101010101010101101;
#1 $display("%b", po);
# 1  pi=24'b001101001101110110100001;
#1 $display("%b", po);
# 1  pi=24'b110011100001100111110100;
#1 $display("%b", po);
# 1  pi=24'b001100111100101001100011;
#1 $display("%b", po);
# 1  pi=24'b000100101101001111111101;
#1 $display("%b", po);
# 1  pi=24'b110111101000011010100011;
#1 $display("%b", po);
# 1  pi=24'b000010001101101111101101;
#1 $display("%b", po);
# 1  pi=24'b111000101101101100110001;
#1 $display("%b", po);
# 1  pi=24'b010101101000011110011001;
#1 $display("%b", po);
# 1  pi=24'b011000001010110010000111;
#1 $display("%b", po);
# 1  pi=24'b111101110111101001111111;
#1 $display("%b", po);
# 1  pi=24'b101101111001011101111101;
#1 $display("%b", po);
# 1  pi=24'b010011110011111001101011;
#1 $display("%b", po);
# 1  pi=24'b011101101010101010001001;
#1 $display("%b", po);
# 1  pi=24'b001001000100101110001100;
#1 $display("%b", po);
# 1  pi=24'b010011110011000110110110;
#1 $display("%b", po);
# 1  pi=24'b110101110000110111011010;
#1 $display("%b", po);
# 1  pi=24'b101100000010101110001000;
#1 $display("%b", po);
# 1  pi=24'b000111000101010000000010;
#1 $display("%b", po);
# 1  pi=24'b011011001100101101001011;
#1 $display("%b", po);
# 1  pi=24'b110111010100111000011100;
#1 $display("%b", po);
# 1  pi=24'b011011100100111100110110;
#1 $display("%b", po);
# 1  pi=24'b000000100010111001100011;
#1 $display("%b", po);
# 1  pi=24'b111101111101111100001011;
#1 $display("%b", po);
# 1  pi=24'b011011011000100110001111;
#1 $display("%b", po);
# 1  pi=24'b110101110110000011011000;
#1 $display("%b", po);
# 1  pi=24'b110101011100000010011011;
#1 $display("%b", po);
# 1  pi=24'b100111001111100110101011;
#1 $display("%b", po);
# 1  pi=24'b110010110110111101011011;
#1 $display("%b", po);
# 1  pi=24'b100010001001001110100100;
#1 $display("%b", po);
# 1  pi=24'b111000110001111110011101;
#1 $display("%b", po);
# 1  pi=24'b101000100011000001100100;
#1 $display("%b", po);
# 1  pi=24'b101011110011100001000101;
#1 $display("%b", po);
# 1  pi=24'b000001000010111010001010;
#1 $display("%b", po);
# 1  pi=24'b001100010101100010110111;
#1 $display("%b", po);
# 1  pi=24'b101011100111111001101000;
#1 $display("%b", po);
# 1  pi=24'b101100011000101011111000;
#1 $display("%b", po);
# 1  pi=24'b110110010000101010110010;
#1 $display("%b", po);
# 1  pi=24'b000011100100010001001010;
#1 $display("%b", po);
# 1  pi=24'b011001111111101100011101;
#1 $display("%b", po);
# 1  pi=24'b111011000110001000010111;
#1 $display("%b", po);
# 1  pi=24'b110001000001101011101110;
#1 $display("%b", po);
# 1  pi=24'b010011000001000011100101;
#1 $display("%b", po);
# 1  pi=24'b110101011011011101010100;
#1 $display("%b", po);
# 1  pi=24'b000001101010100101100110;
#1 $display("%b", po);
# 1  pi=24'b111110100001111000110000;
#1 $display("%b", po);
# 1  pi=24'b010000000000110100011011;
#1 $display("%b", po);
# 1  pi=24'b000111111010001000010101;
#1 $display("%b", po);
# 1  pi=24'b011111100110110000011010;
#1 $display("%b", po);
# 1  pi=24'b010101100110011011111111;
#1 $display("%b", po);
# 1  pi=24'b110100111110010011010111;
#1 $display("%b", po);
# 1  pi=24'b000101010100100000000100;
#1 $display("%b", po);
# 1  pi=24'b111001010001110000100001;
#1 $display("%b", po);
# 1  pi=24'b000101100001111001100110;
#1 $display("%b", po);
# 1  pi=24'b000011001010010001101000;
#1 $display("%b", po);
# 1  pi=24'b110011100001011001001110;
#1 $display("%b", po);
# 1  pi=24'b100011010101101011001000;
#1 $display("%b", po);
# 1  pi=24'b011110111100110011100011;
#1 $display("%b", po);
# 1  pi=24'b010010010000100100010000;
#1 $display("%b", po);
# 1  pi=24'b010100010001110010101111;
#1 $display("%b", po);
# 1  pi=24'b111010101110001011011110;
#1 $display("%b", po);
# 1  pi=24'b111000000011111100111011;
#1 $display("%b", po);
# 1  pi=24'b101100111010000101011001;
#1 $display("%b", po);
# 1  pi=24'b110100111001100000100101;
#1 $display("%b", po);
# 1  pi=24'b101010110111000010000000;
#1 $display("%b", po);
# 1  pi=24'b111100001101101001010110;
#1 $display("%b", po);
# 1  pi=24'b100110100100011000101111;
#1 $display("%b", po);
# 1  pi=24'b000011111000100110010111;
#1 $display("%b", po);
# 1  pi=24'b011011001010100101010101;
#1 $display("%b", po);
# 1  pi=24'b101101010111000101001001;
#1 $display("%b", po);
# 1  pi=24'b011101000110000010000000;
#1 $display("%b", po);
# 1  pi=24'b001110100110011100011101;
#1 $display("%b", po);
# 1  pi=24'b000101101000011110110101;
#1 $display("%b", po);
# 1  pi=24'b111000111001111001111100;
#1 $display("%b", po);
# 1  pi=24'b001111110010000101000101;
#1 $display("%b", po);
# 1  pi=24'b111100101011010111111101;
#1 $display("%b", po);
# 1  pi=24'b100001101000001100011111;
#1 $display("%b", po);
# 1  pi=24'b011101100000100010100011;
#1 $display("%b", po);
# 1  pi=24'b101000011000011101000111;
#1 $display("%b", po);
# 1  pi=24'b001010100000110111101110;
#1 $display("%b", po);
# 1  pi=24'b000011011101000000010111;
#1 $display("%b", po);
# 1  pi=24'b111101010100111110101001;
#1 $display("%b", po);
# 1  pi=24'b011111101011110111100010;
#1 $display("%b", po);
# 1  pi=24'b100000000011101101001010;
#1 $display("%b", po);
# 1  pi=24'b110110010111111000110100;
#1 $display("%b", po);
# 1  pi=24'b111110101101000101100101;
#1 $display("%b", po);
# 1  pi=24'b010010000011110000100111;
#1 $display("%b", po);
# 1  pi=24'b101000100100001101101100;
#1 $display("%b", po);
# 1  pi=24'b001000110111011110101011;
#1 $display("%b", po);
# 1  pi=24'b100110101101001001000011;
#1 $display("%b", po);
# 1  pi=24'b011011001001101101101000;
#1 $display("%b", po);
# 1  pi=24'b101101111111001100010010;
#1 $display("%b", po);
# 1  pi=24'b010111000011010101101001;
#1 $display("%b", po);
# 1  pi=24'b001100010010011001001000;
#1 $display("%b", po);
# 1  pi=24'b010101111011011001011111;
#1 $display("%b", po);
# 1  pi=24'b010011101110111100001001;
#1 $display("%b", po);
# 1  pi=24'b100111011000110000011011;
#1 $display("%b", po);
# 1  pi=24'b001000101100101111110010;
#1 $display("%b", po);
# 1  pi=24'b101001110001100001011001;
#1 $display("%b", po);
# 1  pi=24'b111000011111010100000111;
#1 $display("%b", po);
# 1  pi=24'b011001000011011010111000;
#1 $display("%b", po);
# 1  pi=24'b111010110101010101111110;
#1 $display("%b", po);
# 1  pi=24'b001010001111011101001101;
#1 $display("%b", po);
# 1  pi=24'b000111000010110101110011;
#1 $display("%b", po);
# 1  pi=24'b001001010010111001101111;
#1 $display("%b", po);
# 1  pi=24'b100101111110011100001001;
#1 $display("%b", po);
# 1  pi=24'b000111100110101000100010;
#1 $display("%b", po);
# 1  pi=24'b011111100010001001011100;
#1 $display("%b", po);
# 1  pi=24'b110000101011001011001111;
#1 $display("%b", po);
# 1  pi=24'b101001010110101101111000;
#1 $display("%b", po);
# 1  pi=24'b101101011111001001110000;
#1 $display("%b", po);
# 1  pi=24'b111111111100000001110100;
#1 $display("%b", po);
# 1  pi=24'b001111100000011100100101;
#1 $display("%b", po);
# 1  pi=24'b010100100110001010000011;
#1 $display("%b", po);
# 1  pi=24'b000010100111011000101110;
#1 $display("%b", po);
# 1  pi=24'b011101101011011001000000;
#1 $display("%b", po);
# 1  pi=24'b001000001100101010110001;
#1 $display("%b", po);
# 1  pi=24'b001110100001000010010011;
#1 $display("%b", po);
# 1  pi=24'b011000100110111100101101;
#1 $display("%b", po);
# 1  pi=24'b000110001100000111001100;
#1 $display("%b", po);
# 1  pi=24'b001101010110100111110101;
#1 $display("%b", po);
# 1  pi=24'b010000001010010101011011;
#1 $display("%b", po);
# 1  pi=24'b101000110110000001111111;
#1 $display("%b", po);
# 1  pi=24'b100100110010000011100110;
#1 $display("%b", po);
# 1  pi=24'b101000100100100011000110;
#1 $display("%b", po);
# 1  pi=24'b100111001010111110100011;
#1 $display("%b", po);
# 1  pi=24'b110000101001101111100011;
#1 $display("%b", po);
# 1  pi=24'b000000001011000100111101;
#1 $display("%b", po);
# 1  pi=24'b011000010010101011010011;
#1 $display("%b", po);
# 1  pi=24'b010101110011101011101011;
#1 $display("%b", po);
# 1  pi=24'b001100111111101000000100;
#1 $display("%b", po);
# 1  pi=24'b100101000001110011010000;
#1 $display("%b", po);
# 1  pi=24'b011111010011101001001001;
#1 $display("%b", po);
# 1  pi=24'b100010111111011111000000;
#1 $display("%b", po);
# 1  pi=24'b010001010101011010000110;
#1 $display("%b", po);
# 1  pi=24'b000010101001101110100000;
#1 $display("%b", po);
# 1  pi=24'b110110010100111110010100;
#1 $display("%b", po);
# 1  pi=24'b111001101111010110100000;
#1 $display("%b", po);
# 1  pi=24'b110110000001110001100100;
#1 $display("%b", po);
# 1  pi=24'b101110111111011001101000;
#1 $display("%b", po);
# 1  pi=24'b001101000101010111100001;
#1 $display("%b", po);
# 1  pi=24'b011001000000101010001001;
#1 $display("%b", po);
# 1  pi=24'b101001010001001011101110;
#1 $display("%b", po);
# 1  pi=24'b100110111010000010011110;
#1 $display("%b", po);
# 1  pi=24'b100101001110010000011100;
#1 $display("%b", po);
# 1  pi=24'b001101011011011101001001;
#1 $display("%b", po);
# 1  pi=24'b001000110001100111010110;
#1 $display("%b", po);
# 1  pi=24'b011011100001100010101101;
#1 $display("%b", po);
end
endmodule
